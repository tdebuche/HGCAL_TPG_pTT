parameter integer matrixE [0:1725] = {
/* num inputs = 96(in0-in95) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 3 */
//* total number of input in adders 622 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	2,28,3,47,1,
/* out0003_em-eta3-phi0*/	3,27,1,28,2,47,7,
/* out0004_em-eta4-phi0*/	3,27,3,46,12,47,8,
/* out0005_em-eta5-phi0*/	3,26,2,30,1,46,4,
/* out0006_em-eta6-phi0*/	1,30,11,
/* out0007_em-eta7-phi0*/	3,25,1,29,2,30,3,
/* out0008_em-eta8-phi0*/	1,29,4,
/* out0009_em-eta9-phi0*/	2,2,1,29,3,
/* out0010_em-eta10-phi0*/	1,2,3,
/* out0011_em-eta11-phi0*/	1,2,3,
/* out0012_em-eta12-phi0*/	2,1,1,2,2,
/* out0013_em-eta13-phi0*/	1,1,2,
/* out0014_em-eta14-phi0*/	1,1,2,
/* out0015_em-eta15-phi0*/	1,1,2,
/* out0016_em-eta16-phi0*/	2,0,1,1,1,
/* out0017_em-eta17-phi0*/	1,0,2,
/* out0018_em-eta18-phi0*/	1,0,1,
/* out0019_em-eta19-phi0*/	1,0,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	1,28,7,
/* out0023_em-eta3-phi1*/	3,24,2,27,4,28,4,
/* out0024_em-eta4-phi1*/	2,26,1,27,7,
/* out0025_em-eta5-phi1*/	1,26,7,
/* out0026_em-eta6-phi1*/	3,25,2,26,3,30,1,
/* out0027_em-eta7-phi1*/	1,25,5,
/* out0028_em-eta8-phi1*/	3,6,1,25,2,29,1,
/* out0029_em-eta9-phi1*/	2,6,3,29,6,
/* out0030_em-eta10-phi1*/	2,2,1,6,2,
/* out0031_em-eta11-phi1*/	2,2,5,5,1,
/* out0032_em-eta12-phi1*/	3,1,1,2,1,5,2,
/* out0033_em-eta13-phi1*/	2,1,2,5,1,
/* out0034_em-eta14-phi1*/	1,1,2,
/* out0035_em-eta15-phi1*/	1,1,1,
/* out0036_em-eta16-phi1*/	2,0,1,1,1,
/* out0037_em-eta17-phi1*/	1,0,2,
/* out0038_em-eta18-phi1*/	1,0,1,
/* out0039_em-eta19-phi1*/	1,0,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	2,24,3,34,1,
/* out0043_em-eta3-phi2*/	1,24,10,
/* out0044_em-eta4-phi2*/	2,23,8,27,1,
/* out0045_em-eta5-phi2*/	3,22,2,23,3,26,2,
/* out0046_em-eta6-phi2*/	3,22,4,25,1,26,1,
/* out0047_em-eta7-phi2*/	2,21,1,25,4,
/* out0048_em-eta8-phi2*/	3,6,2,21,1,25,1,
/* out0049_em-eta9-phi2*/	1,6,3,
/* out0050_em-eta10-phi2*/	1,6,2,
/* out0051_em-eta11-phi2*/	1,5,2,
/* out0052_em-eta12-phi2*/	1,5,2,
/* out0053_em-eta13-phi2*/	1,5,2,
/* out0054_em-eta14-phi2*/	2,1,1,4,1,
/* out0055_em-eta15-phi2*/	1,4,1,
/* out0056_em-eta16-phi2*/	1,4,1,
/* out0057_em-eta17-phi2*/	2,0,1,4,1,
/* out0058_em-eta18-phi2*/	1,0,1,
/* out0059_em-eta19-phi2*/	1,0,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	1,34,13,
/* out0063_em-eta3-phi3*/	3,24,1,33,8,34,1,
/* out0064_em-eta4-phi3*/	3,23,4,32,2,33,2,
/* out0065_em-eta5-phi3*/	3,22,4,23,1,32,2,
/* out0066_em-eta6-phi3*/	1,22,5,
/* out0067_em-eta7-phi3*/	1,21,4,
/* out0068_em-eta8-phi3*/	1,21,4,
/* out0069_em-eta9-phi3*/	2,6,2,11,1,
/* out0070_em-eta10-phi3*/	2,6,1,11,2,
/* out0071_em-eta11-phi3*/	1,5,2,
/* out0072_em-eta12-phi3*/	1,5,2,
/* out0073_em-eta13-phi3*/	1,5,1,
/* out0074_em-eta14-phi3*/	1,4,1,
/* out0075_em-eta15-phi3*/	1,4,1,
/* out0076_em-eta16-phi3*/	1,4,1,
/* out0077_em-eta17-phi3*/	1,4,1,
/* out0078_em-eta18-phi3*/	2,0,1,3,1,
/* out0079_em-eta19-phi3*/	1,0,2,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	2,34,1,38,9,
/* out0083_em-eta3-phi4*/	3,33,5,36,3,38,3,
/* out0084_em-eta4-phi4*/	3,32,6,33,1,36,1,
/* out0085_em-eta5-phi4*/	2,31,1,32,5,
/* out0086_em-eta6-phi4*/	2,22,1,31,5,
/* out0087_em-eta7-phi4*/	2,21,3,31,1,
/* out0088_em-eta8-phi4*/	1,21,3,
/* out0089_em-eta9-phi4*/	1,11,3,
/* out0090_em-eta10-phi4*/	1,11,3,
/* out0091_em-eta11-phi4*/	1,11,1,
/* out0092_em-eta12-phi4*/	2,5,1,10,1,
/* out0093_em-eta13-phi4*/	1,10,1,
/* out0094_em-eta14-phi4*/	1,4,1,
/* out0095_em-eta15-phi4*/	1,4,1,
/* out0096_em-eta16-phi4*/	1,4,1,
/* out0097_em-eta17-phi4*/	1,4,1,
/* out0098_em-eta18-phi4*/	1,3,2,
/* out0099_em-eta19-phi4*/	1,3,1,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	2,38,3,39,4,
/* out0103_em-eta3-phi5*/	3,36,8,38,1,39,4,
/* out0104_em-eta4-phi5*/	3,32,1,35,4,36,4,
/* out0105_em-eta5-phi5*/	2,31,2,35,4,
/* out0106_em-eta6-phi5*/	1,31,5,
/* out0107_em-eta7-phi5*/	2,31,2,40,3,
/* out0108_em-eta8-phi5*/	1,40,4,
/* out0109_em-eta9-phi5*/	2,11,2,40,1,
/* out0110_em-eta10-phi5*/	1,11,3,
/* out0111_em-eta11-phi5*/	2,10,2,11,1,
/* out0112_em-eta12-phi5*/	1,10,2,
/* out0113_em-eta13-phi5*/	1,10,1,
/* out0114_em-eta14-phi5*/	2,4,1,10,1,
/* out0115_em-eta15-phi5*/	1,4,1,
/* out0116_em-eta16-phi5*/	1,4,1,
/* out0117_em-eta17-phi5*/	2,3,1,4,1,
/* out0118_em-eta18-phi5*/	1,3,2,
/* out0119_em-eta19-phi5*/	1,3,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	2,39,4,44,3,
/* out0123_em-eta3-phi6*/	3,37,8,39,4,44,1,
/* out0124_em-eta4-phi6*/	3,35,4,37,4,42,1,
/* out0125_em-eta5-phi6*/	2,35,4,41,2,
/* out0126_em-eta6-phi6*/	1,41,5,
/* out0127_em-eta7-phi6*/	2,40,3,41,2,
/* out0128_em-eta8-phi6*/	1,40,4,
/* out0129_em-eta9-phi6*/	2,12,2,40,1,
/* out0130_em-eta10-phi6*/	1,12,3,
/* out0131_em-eta11-phi6*/	2,10,2,12,1,
/* out0132_em-eta12-phi6*/	1,10,2,
/* out0133_em-eta13-phi6*/	1,10,1,
/* out0134_em-eta14-phi6*/	2,7,1,10,1,
/* out0135_em-eta15-phi6*/	1,7,1,
/* out0136_em-eta16-phi6*/	1,7,1,
/* out0137_em-eta17-phi6*/	2,3,1,7,1,
/* out0138_em-eta18-phi6*/	1,3,2,
/* out0139_em-eta19-phi6*/	1,3,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	2,44,9,45,1,
/* out0143_em-eta3-phi7*/	3,37,3,43,5,44,3,
/* out0144_em-eta4-phi7*/	3,37,1,42,6,43,1,
/* out0145_em-eta5-phi7*/	2,41,1,42,5,
/* out0146_em-eta6-phi7*/	2,18,1,41,5,
/* out0147_em-eta7-phi7*/	2,17,3,41,1,
/* out0148_em-eta8-phi7*/	1,17,3,
/* out0149_em-eta9-phi7*/	1,12,3,
/* out0150_em-eta10-phi7*/	1,12,3,
/* out0151_em-eta11-phi7*/	1,12,1,
/* out0152_em-eta12-phi7*/	2,8,1,10,1,
/* out0153_em-eta13-phi7*/	1,10,1,
/* out0154_em-eta14-phi7*/	1,7,1,
/* out0155_em-eta15-phi7*/	1,7,1,
/* out0156_em-eta16-phi7*/	1,7,1,
/* out0157_em-eta17-phi7*/	1,7,1,
/* out0158_em-eta18-phi7*/	1,3,2,
/* out0159_em-eta19-phi7*/	1,3,1,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	1,45,13,
/* out0163_em-eta3-phi8*/	3,20,1,43,8,45,1,
/* out0164_em-eta4-phi8*/	3,19,4,42,2,43,2,
/* out0165_em-eta5-phi8*/	3,18,4,19,1,42,2,
/* out0166_em-eta6-phi8*/	1,18,5,
/* out0167_em-eta7-phi8*/	1,17,4,
/* out0168_em-eta8-phi8*/	1,17,4,
/* out0169_em-eta9-phi8*/	2,9,2,12,1,
/* out0170_em-eta10-phi8*/	2,9,1,12,2,
/* out0171_em-eta11-phi8*/	1,8,2,
/* out0172_em-eta12-phi8*/	1,8,2,
/* out0173_em-eta13-phi8*/	1,8,1,
/* out0174_em-eta14-phi8*/	1,7,1,
/* out0175_em-eta15-phi8*/	1,7,1,
/* out0176_em-eta16-phi8*/	1,7,1,
/* out0177_em-eta17-phi8*/	1,7,1,
/* out0178_em-eta18-phi8*/	1,3,1,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	2,20,3,45,1,
/* out0183_em-eta3-phi9*/	1,20,10,
/* out0184_em-eta4-phi9*/	2,15,1,19,8,
/* out0185_em-eta5-phi9*/	3,14,2,18,2,19,3,
/* out0186_em-eta6-phi9*/	3,13,1,14,1,18,4,
/* out0187_em-eta7-phi9*/	2,13,4,17,1,
/* out0188_em-eta8-phi9*/	3,9,2,13,1,17,1,
/* out0189_em-eta9-phi9*/	1,9,3,
/* out0190_em-eta10-phi9*/	1,9,2,
/* out0191_em-eta11-phi9*/	1,8,2,
/* out0192_em-eta12-phi9*/	1,8,2,
/* out0193_em-eta13-phi9*/	1,8,2,
/* out0194_em-eta14-phi9*/	1,7,1,
/* out0195_em-eta15-phi9*/	1,7,1,
/* out0196_em-eta16-phi9*/	1,7,1,
/* out0197_em-eta17-phi9*/	1,7,1,
/* out0198_em-eta18-phi9*/	1,48,1,
/* out0199_em-eta19-phi9*/	0,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	1,16,3,
/* out0203_em-eta3-phi10*/	3,15,4,16,8,20,2,
/* out0204_em-eta4-phi10*/	2,14,1,15,7,
/* out0205_em-eta5-phi10*/	1,14,7,
/* out0206_em-eta6-phi10*/	2,13,2,14,3,
/* out0207_em-eta7-phi10*/	1,13,5,
/* out0208_em-eta8-phi10*/	3,9,1,13,2,77,1,
/* out0209_em-eta9-phi10*/	1,9,3,
/* out0210_em-eta10-phi10*/	2,9,2,50,1,
/* out0211_em-eta11-phi10*/	2,8,1,50,1,
/* out0212_em-eta12-phi10*/	1,8,2,
/* out0213_em-eta13-phi10*/	2,8,1,49,1,
/* out0214_em-eta14-phi10*/	1,49,1,
/* out0215_em-eta15-phi10*/	1,49,1,
/* out0216_em-eta16-phi10*/	1,48,1,
/* out0217_em-eta17-phi10*/	1,48,1,
/* out0218_em-eta18-phi10*/	1,48,1,
/* out0219_em-eta19-phi10*/	0,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	1,16,1,
/* out0223_em-eta3-phi11*/	3,15,1,16,4,95,7,
/* out0224_em-eta4-phi11*/	3,15,3,94,4,95,1,
/* out0225_em-eta5-phi11*/	3,14,2,78,1,94,4,
/* out0226_em-eta6-phi11*/	1,78,5,
/* out0227_em-eta7-phi11*/	3,13,1,77,1,78,2,
/* out0228_em-eta8-phi11*/	1,77,4,
/* out0229_em-eta9-phi11*/	1,77,2,
/* out0230_em-eta10-phi11*/	1,50,3,
/* out0231_em-eta11-phi11*/	1,50,2,
/* out0232_em-eta12-phi11*/	2,49,1,50,1,
/* out0233_em-eta13-phi11*/	1,49,2,
/* out0234_em-eta14-phi11*/	1,49,1,
/* out0235_em-eta15-phi11*/	1,49,1,
/* out0236_em-eta16-phi11*/	1,48,1,
/* out0237_em-eta17-phi11*/	1,48,1,
/* out0238_em-eta18-phi11*/	1,48,1,
/* out0239_em-eta19-phi11*/	1,48,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	1,76,3,
/* out0243_em-eta3-phi12*/	3,75,1,76,2,95,7,
/* out0244_em-eta4-phi12*/	3,75,3,94,4,95,1,
/* out0245_em-eta5-phi12*/	3,74,2,78,1,94,4,
/* out0246_em-eta6-phi12*/	1,78,5,
/* out0247_em-eta7-phi12*/	3,73,1,77,1,78,2,
/* out0248_em-eta8-phi12*/	1,77,4,
/* out0249_em-eta9-phi12*/	1,77,2,
/* out0250_em-eta10-phi12*/	1,50,3,
/* out0251_em-eta11-phi12*/	1,50,2,
/* out0252_em-eta12-phi12*/	2,49,1,50,1,
/* out0253_em-eta13-phi12*/	1,49,2,
/* out0254_em-eta14-phi12*/	1,49,1,
/* out0255_em-eta15-phi12*/	1,49,1,
/* out0256_em-eta16-phi12*/	1,48,1,
/* out0257_em-eta17-phi12*/	1,48,1,
/* out0258_em-eta18-phi12*/	1,48,1,
/* out0259_em-eta19-phi12*/	1,48,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	1,76,7,
/* out0263_em-eta3-phi13*/	3,72,2,75,4,76,4,
/* out0264_em-eta4-phi13*/	2,74,1,75,7,
/* out0265_em-eta5-phi13*/	1,74,7,
/* out0266_em-eta6-phi13*/	2,73,2,74,3,
/* out0267_em-eta7-phi13*/	1,73,5,
/* out0268_em-eta8-phi13*/	3,54,1,73,2,77,1,
/* out0269_em-eta9-phi13*/	1,54,3,
/* out0270_em-eta10-phi13*/	2,50,1,54,2,
/* out0271_em-eta11-phi13*/	2,50,1,53,1,
/* out0272_em-eta12-phi13*/	1,53,2,
/* out0273_em-eta13-phi13*/	2,49,1,53,1,
/* out0274_em-eta14-phi13*/	1,49,1,
/* out0275_em-eta15-phi13*/	1,49,1,
/* out0276_em-eta16-phi13*/	1,48,1,
/* out0277_em-eta17-phi13*/	1,48,1,
/* out0278_em-eta18-phi13*/	1,48,1,
/* out0279_em-eta19-phi13*/	0,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	2,72,3,82,1,
/* out0283_em-eta3-phi14*/	1,72,10,
/* out0284_em-eta4-phi14*/	2,71,8,75,1,
/* out0285_em-eta5-phi14*/	3,70,2,71,3,74,2,
/* out0286_em-eta6-phi14*/	3,70,4,73,1,74,1,
/* out0287_em-eta7-phi14*/	2,69,1,73,4,
/* out0288_em-eta8-phi14*/	3,54,2,69,1,73,1,
/* out0289_em-eta9-phi14*/	1,54,3,
/* out0290_em-eta10-phi14*/	1,54,2,
/* out0291_em-eta11-phi14*/	1,53,2,
/* out0292_em-eta12-phi14*/	1,53,2,
/* out0293_em-eta13-phi14*/	1,53,2,
/* out0294_em-eta14-phi14*/	1,52,1,
/* out0295_em-eta15-phi14*/	1,52,1,
/* out0296_em-eta16-phi14*/	1,52,1,
/* out0297_em-eta17-phi14*/	1,52,1,
/* out0298_em-eta18-phi14*/	1,48,1,
/* out0299_em-eta19-phi14*/	0,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	1,82,13,
/* out0303_em-eta3-phi15*/	3,72,1,81,8,82,1,
/* out0304_em-eta4-phi15*/	3,71,4,80,2,81,2,
/* out0305_em-eta5-phi15*/	3,70,4,71,1,80,2,
/* out0306_em-eta6-phi15*/	1,70,5,
/* out0307_em-eta7-phi15*/	1,69,4,
/* out0308_em-eta8-phi15*/	1,69,4,
/* out0309_em-eta9-phi15*/	2,54,2,60,1,
/* out0310_em-eta10-phi15*/	2,54,1,60,2,
/* out0311_em-eta11-phi15*/	1,53,2,
/* out0312_em-eta12-phi15*/	1,53,2,
/* out0313_em-eta13-phi15*/	1,53,1,
/* out0314_em-eta14-phi15*/	1,52,1,
/* out0315_em-eta15-phi15*/	1,52,1,
/* out0316_em-eta16-phi15*/	1,52,1,
/* out0317_em-eta17-phi15*/	1,52,1,
/* out0318_em-eta18-phi15*/	1,51,1,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	2,82,1,87,9,
/* out0323_em-eta3-phi16*/	3,81,5,85,3,87,3,
/* out0324_em-eta4-phi16*/	3,80,6,81,1,85,1,
/* out0325_em-eta5-phi16*/	2,79,1,80,5,
/* out0326_em-eta6-phi16*/	2,70,1,79,5,
/* out0327_em-eta7-phi16*/	2,69,3,79,1,
/* out0328_em-eta8-phi16*/	1,69,3,
/* out0329_em-eta9-phi16*/	1,60,3,
/* out0330_em-eta10-phi16*/	1,60,3,
/* out0331_em-eta11-phi16*/	1,60,1,
/* out0332_em-eta12-phi16*/	2,53,1,58,1,
/* out0333_em-eta13-phi16*/	1,58,1,
/* out0334_em-eta14-phi16*/	1,52,1,
/* out0335_em-eta15-phi16*/	1,52,1,
/* out0336_em-eta16-phi16*/	1,52,1,
/* out0337_em-eta17-phi16*/	1,52,1,
/* out0338_em-eta18-phi16*/	1,51,2,
/* out0339_em-eta19-phi16*/	1,51,1,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	2,86,4,87,3,
/* out0343_em-eta3-phi17*/	3,85,8,86,4,87,1,
/* out0344_em-eta4-phi17*/	3,80,1,83,4,85,4,
/* out0345_em-eta5-phi17*/	2,79,2,83,4,
/* out0346_em-eta6-phi17*/	1,79,5,
/* out0347_em-eta7-phi17*/	2,79,2,88,3,
/* out0348_em-eta8-phi17*/	1,88,4,
/* out0349_em-eta9-phi17*/	2,60,2,88,1,
/* out0350_em-eta10-phi17*/	1,60,3,
/* out0351_em-eta11-phi17*/	2,58,2,60,1,
/* out0352_em-eta12-phi17*/	1,58,2,
/* out0353_em-eta13-phi17*/	1,58,1,
/* out0354_em-eta14-phi17*/	2,52,1,58,1,
/* out0355_em-eta15-phi17*/	1,52,1,
/* out0356_em-eta16-phi17*/	1,52,1,
/* out0357_em-eta17-phi17*/	2,51,1,52,1,
/* out0358_em-eta18-phi17*/	1,51,2,
/* out0359_em-eta19-phi17*/	1,51,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	2,86,4,93,3,
/* out0363_em-eta3-phi18*/	3,84,8,86,4,93,1,
/* out0364_em-eta4-phi18*/	3,83,4,84,4,90,1,
/* out0365_em-eta5-phi18*/	2,83,4,89,2,
/* out0366_em-eta6-phi18*/	1,89,5,
/* out0367_em-eta7-phi18*/	2,88,3,89,2,
/* out0368_em-eta8-phi18*/	1,88,4,
/* out0369_em-eta9-phi18*/	2,59,2,88,1,
/* out0370_em-eta10-phi18*/	1,59,3,
/* out0371_em-eta11-phi18*/	2,58,2,59,1,
/* out0372_em-eta12-phi18*/	1,58,2,
/* out0373_em-eta13-phi18*/	1,58,1,
/* out0374_em-eta14-phi18*/	2,55,1,58,1,
/* out0375_em-eta15-phi18*/	1,55,1,
/* out0376_em-eta16-phi18*/	1,55,1,
/* out0377_em-eta17-phi18*/	2,51,1,55,1,
/* out0378_em-eta18-phi18*/	1,51,2,
/* out0379_em-eta19-phi18*/	1,51,1,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	2,92,1,93,9,
/* out0383_em-eta3-phi19*/	3,84,3,91,5,93,3,
/* out0384_em-eta4-phi19*/	3,84,1,90,6,91,1,
/* out0385_em-eta5-phi19*/	2,89,1,90,5,
/* out0386_em-eta6-phi19*/	2,66,1,89,5,
/* out0387_em-eta7-phi19*/	2,65,3,89,1,
/* out0388_em-eta8-phi19*/	1,65,3,
/* out0389_em-eta9-phi19*/	1,59,3,
/* out0390_em-eta10-phi19*/	1,59,3,
/* out0391_em-eta11-phi19*/	1,59,1,
/* out0392_em-eta12-phi19*/	2,56,1,58,1,
/* out0393_em-eta13-phi19*/	1,58,1,
/* out0394_em-eta14-phi19*/	1,55,1,
/* out0395_em-eta15-phi19*/	1,55,1,
/* out0396_em-eta16-phi19*/	1,55,1,
/* out0397_em-eta17-phi19*/	1,55,1,
/* out0398_em-eta18-phi19*/	1,51,2,
/* out0399_em-eta19-phi19*/	1,51,1,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	1,92,13,
/* out0403_em-eta3-phi20*/	3,68,1,91,8,92,1,
/* out0404_em-eta4-phi20*/	3,67,4,90,2,91,2,
/* out0405_em-eta5-phi20*/	3,66,4,67,1,90,2,
/* out0406_em-eta6-phi20*/	1,66,5,
/* out0407_em-eta7-phi20*/	1,65,4,
/* out0408_em-eta8-phi20*/	1,65,4,
/* out0409_em-eta9-phi20*/	2,57,2,59,1,
/* out0410_em-eta10-phi20*/	2,57,1,59,2,
/* out0411_em-eta11-phi20*/	1,56,2,
/* out0412_em-eta12-phi20*/	1,56,2,
/* out0413_em-eta13-phi20*/	1,56,1,
/* out0414_em-eta14-phi20*/	1,55,1,
/* out0415_em-eta15-phi20*/	1,55,1,
/* out0416_em-eta16-phi20*/	1,55,1,
/* out0417_em-eta17-phi20*/	1,55,1,
/* out0418_em-eta18-phi20*/	1,51,1,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	2,68,3,92,1,
/* out0423_em-eta3-phi21*/	1,68,10,
/* out0424_em-eta4-phi21*/	2,63,1,67,8,
/* out0425_em-eta5-phi21*/	3,62,2,66,2,67,3,
/* out0426_em-eta6-phi21*/	3,61,1,62,1,66,4,
/* out0427_em-eta7-phi21*/	2,61,4,65,1,
/* out0428_em-eta8-phi21*/	3,57,2,61,1,65,1,
/* out0429_em-eta9-phi21*/	1,57,3,
/* out0430_em-eta10-phi21*/	1,57,2,
/* out0431_em-eta11-phi21*/	1,56,2,
/* out0432_em-eta12-phi21*/	1,56,2,
/* out0433_em-eta13-phi21*/	1,56,2,
/* out0434_em-eta14-phi21*/	1,55,1,
/* out0435_em-eta15-phi21*/	1,55,1,
/* out0436_em-eta16-phi21*/	1,55,1,
/* out0437_em-eta17-phi21*/	1,55,1,
/* out0438_em-eta18-phi21*/	0,
/* out0439_em-eta19-phi21*/	0,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	1,64,3,
/* out0443_em-eta3-phi22*/	3,63,4,64,8,68,2,
/* out0444_em-eta4-phi22*/	2,62,1,63,7,
/* out0445_em-eta5-phi22*/	1,62,7,
/* out0446_em-eta6-phi22*/	2,61,2,62,3,
/* out0447_em-eta7-phi22*/	1,61,5,
/* out0448_em-eta8-phi22*/	2,57,1,61,2,
/* out0449_em-eta9-phi22*/	1,57,3,
/* out0450_em-eta10-phi22*/	1,57,2,
/* out0451_em-eta11-phi22*/	1,56,1,
/* out0452_em-eta12-phi22*/	1,56,2,
/* out0453_em-eta13-phi22*/	1,56,1,
/* out0454_em-eta14-phi22*/	0,
/* out0455_em-eta15-phi22*/	0,
/* out0456_em-eta16-phi22*/	0,
/* out0457_em-eta17-phi22*/	0,
/* out0458_em-eta18-phi22*/	0,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	1,64,1,
/* out0463_em-eta3-phi23*/	2,63,1,64,4,
/* out0464_em-eta4-phi23*/	1,63,3,
/* out0465_em-eta5-phi23*/	1,62,2,
/* out0466_em-eta6-phi23*/	0,
/* out0467_em-eta7-phi23*/	1,61,1,
/* out0468_em-eta8-phi23*/	0,
/* out0469_em-eta9-phi23*/	0,
/* out0470_em-eta10-phi23*/	0,
/* out0471_em-eta11-phi23*/	0,
/* out0472_em-eta12-phi23*/	0,
/* out0473_em-eta13-phi23*/	0,
/* out0474_em-eta14-phi23*/	0,
/* out0475_em-eta15-phi23*/	0,
/* out0476_em-eta16-phi23*/	0,
/* out0477_em-eta17-phi23*/	0,
/* out0478_em-eta18-phi23*/	0,
/* out0479_em-eta19-phi23*/	0
};