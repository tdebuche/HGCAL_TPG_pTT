parameter integer matrixH [0:2340] = {
/* num inputs = 152(in0-in151) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 6 */
//* total number of input in adders 930 */

/* out0000_had-eta0-phi0*/	1, 107, 2, 
/* out0001_had-eta1-phi0*/	2, 106, 2, 107, 6, 
/* out0002_had-eta2-phi0*/	1, 106, 4, 
/* out0003_had-eta3-phi0*/	2, 105, 3, 106, 2, 
/* out0004_had-eta4-phi0*/	1, 105, 4, 
/* out0005_had-eta5-phi0*/	2, 104, 4, 105, 1, 
/* out0006_had-eta6-phi0*/	1, 104, 4, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	2, 47, 8, 99, 8, 
/* out0010_had-eta10-phi0*/	3, 46, 2, 47, 5, 98, 4, 
/* out0011_had-eta11-phi0*/	2, 46, 5, 98, 3, 
/* out0012_had-eta12-phi0*/	3, 45, 1, 46, 4, 97, 3, 
/* out0013_had-eta13-phi0*/	2, 45, 4, 97, 2, 
/* out0014_had-eta14-phi0*/	2, 45, 3, 96, 1, 
/* out0015_had-eta15-phi0*/	3, 44, 2, 45, 1, 96, 2, 
/* out0016_had-eta16-phi0*/	2, 44, 2, 96, 1, 
/* out0017_had-eta17-phi0*/	2, 44, 2, 95, 1, 
/* out0018_had-eta18-phi0*/	2, 44, 1, 95, 2, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	1, 107, 2, 
/* out0021_had-eta1-phi1*/	2, 106, 2, 107, 6, 
/* out0022_had-eta2-phi1*/	1, 106, 4, 
/* out0023_had-eta3-phi1*/	2, 105, 3, 106, 2, 
/* out0024_had-eta4-phi1*/	1, 105, 4, 
/* out0025_had-eta5-phi1*/	2, 104, 4, 105, 1, 
/* out0026_had-eta6-phi1*/	1, 104, 4, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	1, 43, 1, 
/* out0029_had-eta9-phi1*/	5, 42, 1, 43, 8, 47, 2, 93, 2, 99, 8, 
/* out0030_had-eta10-phi1*/	4, 42, 4, 47, 1, 93, 1, 98, 5, 
/* out0031_had-eta11-phi1*/	5, 41, 1, 42, 1, 46, 3, 97, 1, 98, 4, 
/* out0032_had-eta12-phi1*/	4, 41, 2, 45, 1, 46, 2, 97, 4, 
/* out0033_had-eta13-phi1*/	2, 45, 3, 97, 3, 
/* out0034_had-eta14-phi1*/	2, 45, 3, 96, 3, 
/* out0035_had-eta15-phi1*/	2, 44, 2, 96, 2, 
/* out0036_had-eta16-phi1*/	2, 44, 2, 96, 2, 
/* out0037_had-eta17-phi1*/	2, 44, 2, 95, 3, 
/* out0038_had-eta18-phi1*/	2, 44, 1, 95, 2, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	1, 111, 2, 
/* out0041_had-eta1-phi2*/	2, 110, 2, 111, 6, 
/* out0042_had-eta2-phi2*/	1, 110, 4, 
/* out0043_had-eta3-phi2*/	2, 109, 3, 110, 2, 
/* out0044_had-eta4-phi2*/	1, 109, 4, 
/* out0045_had-eta5-phi2*/	2, 108, 4, 109, 1, 
/* out0046_had-eta6-phi2*/	1, 108, 4, 
/* out0047_had-eta7-phi2*/	0, 
/* out0048_had-eta8-phi2*/	2, 37, 1, 43, 2, 
/* out0049_had-eta9-phi2*/	4, 37, 3, 42, 2, 43, 5, 93, 6, 
/* out0050_had-eta10-phi2*/	3, 42, 5, 91, 2, 93, 4, 
/* out0051_had-eta11-phi2*/	3, 41, 2, 42, 2, 91, 5, 
/* out0052_had-eta12-phi2*/	4, 41, 4, 90, 1, 91, 2, 97, 2, 
/* out0053_had-eta13-phi2*/	4, 40, 1, 41, 2, 90, 2, 97, 1, 
/* out0054_had-eta14-phi2*/	3, 40, 3, 90, 1, 96, 2, 
/* out0055_had-eta15-phi2*/	2, 40, 2, 96, 2, 
/* out0056_had-eta16-phi2*/	3, 44, 1, 95, 1, 96, 1, 
/* out0057_had-eta17-phi2*/	3, 39, 1, 44, 1, 95, 3, 
/* out0058_had-eta18-phi2*/	2, 39, 1, 95, 1, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	1, 111, 2, 
/* out0061_had-eta1-phi3*/	2, 110, 2, 111, 6, 
/* out0062_had-eta2-phi3*/	1, 110, 4, 
/* out0063_had-eta3-phi3*/	2, 109, 3, 110, 2, 
/* out0064_had-eta4-phi3*/	1, 109, 4, 
/* out0065_had-eta5-phi3*/	2, 108, 4, 109, 1, 
/* out0066_had-eta6-phi3*/	1, 108, 4, 
/* out0067_had-eta7-phi3*/	0, 
/* out0068_had-eta8-phi3*/	1, 37, 1, 
/* out0069_had-eta9-phi3*/	3, 37, 8, 93, 2, 94, 2, 
/* out0070_had-eta10-phi3*/	6, 36, 4, 37, 1, 42, 1, 91, 1, 93, 1, 94, 4, 
/* out0071_had-eta11-phi3*/	3, 36, 4, 41, 1, 91, 4, 
/* out0072_had-eta12-phi3*/	4, 35, 1, 41, 3, 90, 2, 91, 2, 
/* out0073_had-eta13-phi3*/	4, 35, 1, 40, 1, 41, 1, 90, 3, 
/* out0074_had-eta14-phi3*/	2, 40, 3, 90, 2, 
/* out0075_had-eta15-phi3*/	2, 40, 2, 89, 2, 
/* out0076_had-eta16-phi3*/	3, 39, 2, 40, 1, 89, 2, 
/* out0077_had-eta17-phi3*/	3, 39, 2, 89, 1, 95, 2, 
/* out0078_had-eta18-phi3*/	2, 39, 1, 95, 1, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	1, 115, 2, 
/* out0081_had-eta1-phi4*/	2, 114, 2, 115, 6, 
/* out0082_had-eta2-phi4*/	1, 114, 4, 
/* out0083_had-eta3-phi4*/	2, 113, 3, 114, 2, 
/* out0084_had-eta4-phi4*/	1, 113, 4, 
/* out0085_had-eta5-phi4*/	2, 112, 4, 113, 1, 
/* out0086_had-eta6-phi4*/	1, 112, 4, 
/* out0087_had-eta7-phi4*/	0, 
/* out0088_had-eta8-phi4*/	0, 
/* out0089_had-eta9-phi4*/	3, 37, 2, 38, 5, 94, 4, 
/* out0090_had-eta10-phi4*/	3, 36, 4, 38, 2, 94, 6, 
/* out0091_had-eta11-phi4*/	3, 35, 1, 36, 4, 92, 5, 
/* out0092_had-eta12-phi4*/	3, 35, 4, 90, 1, 92, 4, 
/* out0093_had-eta13-phi4*/	2, 35, 3, 90, 3, 
/* out0094_had-eta14-phi4*/	4, 29, 1, 40, 2, 89, 1, 90, 1, 
/* out0095_had-eta15-phi4*/	3, 29, 1, 40, 1, 89, 2, 
/* out0096_had-eta16-phi4*/	2, 39, 2, 89, 2, 
/* out0097_had-eta17-phi4*/	2, 39, 2, 89, 1, 
/* out0098_had-eta18-phi4*/	1, 39, 1, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	1, 115, 2, 
/* out0101_had-eta1-phi5*/	2, 114, 2, 115, 6, 
/* out0102_had-eta2-phi5*/	1, 114, 4, 
/* out0103_had-eta3-phi5*/	2, 113, 3, 114, 2, 
/* out0104_had-eta4-phi5*/	1, 113, 4, 
/* out0105_had-eta5-phi5*/	2, 112, 4, 113, 1, 
/* out0106_had-eta6-phi5*/	1, 112, 4, 
/* out0107_had-eta7-phi5*/	0, 
/* out0108_had-eta8-phi5*/	0, 
/* out0109_had-eta9-phi5*/	2, 38, 7, 102, 2, 
/* out0110_had-eta10-phi5*/	3, 31, 3, 38, 2, 102, 5, 
/* out0111_had-eta11-phi5*/	3, 31, 4, 92, 4, 102, 1, 
/* out0112_had-eta12-phi5*/	4, 31, 1, 35, 3, 92, 3, 100, 1, 
/* out0113_had-eta13-phi5*/	2, 35, 3, 100, 3, 
/* out0114_had-eta14-phi5*/	2, 29, 3, 100, 3, 
/* out0115_had-eta15-phi5*/	2, 29, 2, 89, 2, 
/* out0116_had-eta16-phi5*/	3, 29, 1, 39, 1, 89, 2, 
/* out0117_had-eta17-phi5*/	2, 39, 2, 89, 1, 
/* out0118_had-eta18-phi5*/	1, 39, 1, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	1, 119, 2, 
/* out0121_had-eta1-phi6*/	2, 118, 2, 119, 6, 
/* out0122_had-eta2-phi6*/	1, 118, 4, 
/* out0123_had-eta3-phi6*/	2, 117, 3, 118, 2, 
/* out0124_had-eta4-phi6*/	1, 117, 4, 
/* out0125_had-eta5-phi6*/	2, 116, 4, 117, 1, 
/* out0126_had-eta6-phi6*/	1, 116, 4, 
/* out0127_had-eta7-phi6*/	0, 
/* out0128_had-eta8-phi6*/	0, 
/* out0129_had-eta9-phi6*/	2, 33, 7, 102, 2, 
/* out0130_had-eta10-phi6*/	3, 31, 3, 33, 2, 102, 5, 
/* out0131_had-eta11-phi6*/	3, 31, 4, 101, 4, 102, 1, 
/* out0132_had-eta12-phi6*/	4, 30, 3, 31, 1, 100, 1, 101, 3, 
/* out0133_had-eta13-phi6*/	2, 30, 3, 100, 3, 
/* out0134_had-eta14-phi6*/	2, 29, 3, 100, 3, 
/* out0135_had-eta15-phi6*/	2, 29, 2, 85, 2, 
/* out0136_had-eta16-phi6*/	3, 24, 1, 29, 1, 85, 2, 
/* out0137_had-eta17-phi6*/	2, 24, 2, 85, 1, 
/* out0138_had-eta18-phi6*/	1, 24, 1, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	1, 119, 2, 
/* out0141_had-eta1-phi7*/	2, 118, 2, 119, 6, 
/* out0142_had-eta2-phi7*/	1, 118, 4, 
/* out0143_had-eta3-phi7*/	2, 117, 3, 118, 2, 
/* out0144_had-eta4-phi7*/	1, 117, 4, 
/* out0145_had-eta5-phi7*/	2, 116, 4, 117, 1, 
/* out0146_had-eta6-phi7*/	1, 116, 4, 
/* out0147_had-eta7-phi7*/	0, 
/* out0148_had-eta8-phi7*/	0, 
/* out0149_had-eta9-phi7*/	3, 33, 5, 34, 2, 103, 4, 
/* out0150_had-eta10-phi7*/	3, 32, 4, 33, 2, 103, 6, 
/* out0151_had-eta11-phi7*/	3, 30, 1, 32, 4, 101, 5, 
/* out0152_had-eta12-phi7*/	3, 30, 4, 86, 1, 101, 4, 
/* out0153_had-eta13-phi7*/	3, 30, 3, 86, 3, 100, 1, 
/* out0154_had-eta14-phi7*/	5, 25, 2, 29, 1, 85, 1, 86, 1, 100, 1, 
/* out0155_had-eta15-phi7*/	3, 25, 1, 29, 1, 85, 2, 
/* out0156_had-eta16-phi7*/	2, 24, 2, 85, 2, 
/* out0157_had-eta17-phi7*/	2, 24, 2, 85, 1, 
/* out0158_had-eta18-phi7*/	1, 24, 1, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	1, 123, 2, 
/* out0161_had-eta1-phi8*/	2, 122, 2, 123, 6, 
/* out0162_had-eta2-phi8*/	1, 122, 4, 
/* out0163_had-eta3-phi8*/	2, 121, 3, 122, 2, 
/* out0164_had-eta4-phi8*/	1, 121, 4, 
/* out0165_had-eta5-phi8*/	2, 120, 4, 121, 1, 
/* out0166_had-eta6-phi8*/	1, 120, 4, 
/* out0167_had-eta7-phi8*/	0, 
/* out0168_had-eta8-phi8*/	1, 34, 1, 
/* out0169_had-eta9-phi8*/	3, 34, 8, 88, 2, 103, 2, 
/* out0170_had-eta10-phi8*/	6, 27, 1, 32, 4, 34, 1, 87, 1, 88, 1, 103, 4, 
/* out0171_had-eta11-phi8*/	3, 26, 1, 32, 4, 87, 4, 
/* out0172_had-eta12-phi8*/	4, 26, 3, 30, 1, 86, 2, 87, 2, 
/* out0173_had-eta13-phi8*/	4, 25, 1, 26, 1, 30, 1, 86, 3, 
/* out0174_had-eta14-phi8*/	2, 25, 3, 86, 2, 
/* out0175_had-eta15-phi8*/	2, 25, 2, 85, 2, 
/* out0176_had-eta16-phi8*/	3, 24, 2, 25, 1, 85, 2, 
/* out0177_had-eta17-phi8*/	3, 24, 2, 80, 2, 85, 1, 
/* out0178_had-eta18-phi8*/	2, 24, 1, 80, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	1, 123, 2, 
/* out0181_had-eta1-phi9*/	2, 122, 2, 123, 6, 
/* out0182_had-eta2-phi9*/	1, 122, 4, 
/* out0183_had-eta3-phi9*/	2, 121, 3, 122, 2, 
/* out0184_had-eta4-phi9*/	1, 121, 4, 
/* out0185_had-eta5-phi9*/	2, 120, 4, 121, 1, 
/* out0186_had-eta6-phi9*/	1, 120, 4, 
/* out0187_had-eta7-phi9*/	0, 
/* out0188_had-eta8-phi9*/	2, 28, 2, 34, 1, 
/* out0189_had-eta9-phi9*/	4, 27, 2, 28, 5, 34, 3, 88, 7, 
/* out0190_had-eta10-phi9*/	3, 27, 5, 87, 2, 88, 4, 
/* out0191_had-eta11-phi9*/	3, 26, 2, 27, 2, 87, 5, 
/* out0192_had-eta12-phi9*/	4, 26, 4, 82, 2, 86, 1, 87, 2, 
/* out0193_had-eta13-phi9*/	4, 25, 1, 26, 2, 82, 1, 86, 2, 
/* out0194_had-eta14-phi9*/	3, 25, 3, 81, 2, 86, 1, 
/* out0195_had-eta15-phi9*/	2, 25, 2, 81, 2, 
/* out0196_had-eta16-phi9*/	3, 20, 1, 80, 1, 81, 1, 
/* out0197_had-eta17-phi9*/	3, 20, 1, 24, 1, 80, 3, 
/* out0198_had-eta18-phi9*/	2, 24, 1, 80, 1, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	1, 127, 2, 
/* out0201_had-eta1-phi10*/	2, 126, 2, 127, 6, 
/* out0202_had-eta2-phi10*/	1, 126, 4, 
/* out0203_had-eta3-phi10*/	2, 125, 3, 126, 2, 
/* out0204_had-eta4-phi10*/	1, 125, 4, 
/* out0205_had-eta5-phi10*/	2, 124, 4, 125, 1, 
/* out0206_had-eta6-phi10*/	1, 124, 4, 
/* out0207_had-eta7-phi10*/	0, 
/* out0208_had-eta8-phi10*/	1, 28, 1, 
/* out0209_had-eta9-phi10*/	5, 23, 2, 27, 1, 28, 8, 84, 8, 88, 2, 
/* out0210_had-eta10-phi10*/	3, 23, 1, 27, 4, 83, 5, 
/* out0211_had-eta11-phi10*/	5, 22, 3, 26, 1, 27, 1, 82, 1, 83, 4, 
/* out0212_had-eta12-phi10*/	4, 21, 1, 22, 1, 26, 2, 82, 4, 
/* out0213_had-eta13-phi10*/	2, 21, 3, 82, 3, 
/* out0214_had-eta14-phi10*/	2, 21, 2, 81, 3, 
/* out0215_had-eta15-phi10*/	2, 20, 2, 81, 2, 
/* out0216_had-eta16-phi10*/	2, 20, 2, 81, 2, 
/* out0217_had-eta17-phi10*/	2, 20, 1, 80, 3, 
/* out0218_had-eta18-phi10*/	2, 20, 1, 80, 2, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	1, 127, 2, 
/* out0221_had-eta1-phi11*/	2, 126, 2, 127, 6, 
/* out0222_had-eta2-phi11*/	1, 126, 4, 
/* out0223_had-eta3-phi11*/	2, 125, 3, 126, 2, 
/* out0224_had-eta4-phi11*/	1, 125, 4, 
/* out0225_had-eta5-phi11*/	2, 124, 4, 125, 1, 
/* out0226_had-eta6-phi11*/	1, 124, 4, 
/* out0227_had-eta7-phi11*/	0, 
/* out0228_had-eta8-phi11*/	0, 
/* out0229_had-eta9-phi11*/	3, 23, 6, 79, 1, 84, 8, 
/* out0230_had-eta10-phi11*/	4, 22, 1, 23, 4, 79, 2, 83, 4, 
/* out0231_had-eta11-phi11*/	3, 22, 5, 78, 1, 83, 3, 
/* out0232_had-eta12-phi11*/	4, 21, 1, 22, 3, 78, 1, 82, 3, 
/* out0233_had-eta13-phi11*/	3, 21, 3, 77, 1, 82, 2, 
/* out0234_had-eta14-phi11*/	3, 21, 3, 77, 1, 81, 1, 
/* out0235_had-eta15-phi11*/	3, 20, 2, 21, 1, 81, 2, 
/* out0236_had-eta16-phi11*/	3, 20, 2, 76, 1, 81, 1, 
/* out0237_had-eta17-phi11*/	3, 20, 1, 76, 1, 80, 1, 
/* out0238_had-eta18-phi11*/	2, 20, 1, 80, 2, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	1, 131, 2, 
/* out0241_had-eta1-phi12*/	2, 130, 2, 131, 6, 
/* out0242_had-eta2-phi12*/	1, 130, 4, 
/* out0243_had-eta3-phi12*/	2, 129, 3, 130, 2, 
/* out0244_had-eta4-phi12*/	1, 129, 4, 
/* out0245_had-eta5-phi12*/	2, 128, 4, 129, 1, 
/* out0246_had-eta6-phi12*/	1, 128, 4, 
/* out0247_had-eta7-phi12*/	0, 
/* out0248_had-eta8-phi12*/	0, 
/* out0249_had-eta9-phi12*/	4, 18, 1, 19, 8, 23, 2, 79, 5, 
/* out0250_had-eta10-phi12*/	3, 18, 4, 23, 1, 79, 5, 
/* out0251_had-eta11-phi12*/	3, 18, 2, 22, 2, 78, 5, 
/* out0252_had-eta12-phi12*/	3, 17, 3, 22, 1, 78, 4, 
/* out0253_had-eta13-phi12*/	3, 17, 2, 21, 1, 77, 3, 
/* out0254_had-eta14-phi12*/	3, 16, 2, 21, 1, 77, 3, 
/* out0255_had-eta15-phi12*/	3, 16, 2, 76, 1, 77, 1, 
/* out0256_had-eta16-phi12*/	3, 16, 1, 20, 1, 76, 2, 
/* out0257_had-eta17-phi12*/	3, 15, 1, 20, 1, 76, 2, 
/* out0258_had-eta18-phi12*/	2, 15, 1, 76, 1, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	1, 131, 2, 
/* out0261_had-eta1-phi13*/	2, 130, 2, 131, 6, 
/* out0262_had-eta2-phi13*/	1, 130, 4, 
/* out0263_had-eta3-phi13*/	2, 129, 3, 130, 2, 
/* out0264_had-eta4-phi13*/	1, 129, 4, 
/* out0265_had-eta5-phi13*/	2, 128, 4, 129, 1, 
/* out0266_had-eta6-phi13*/	1, 128, 4, 
/* out0267_had-eta7-phi13*/	0, 
/* out0268_had-eta8-phi13*/	1, 19, 1, 
/* out0269_had-eta9-phi13*/	5, 14, 2, 18, 1, 19, 7, 75, 9, 79, 1, 
/* out0270_had-eta10-phi13*/	3, 18, 5, 74, 4, 79, 2, 
/* out0271_had-eta11-phi13*/	4, 17, 1, 18, 3, 74, 2, 78, 3, 
/* out0272_had-eta12-phi13*/	3, 17, 4, 73, 2, 78, 2, 
/* out0273_had-eta13-phi13*/	3, 17, 3, 73, 1, 77, 3, 
/* out0274_had-eta14-phi13*/	2, 16, 3, 77, 3, 
/* out0275_had-eta15-phi13*/	4, 16, 2, 72, 1, 76, 1, 77, 1, 
/* out0276_had-eta16-phi13*/	3, 15, 1, 16, 1, 76, 2, 
/* out0277_had-eta17-phi13*/	2, 15, 3, 76, 2, 
/* out0278_had-eta18-phi13*/	2, 15, 1, 76, 1, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	1, 135, 2, 
/* out0281_had-eta1-phi14*/	2, 134, 2, 135, 6, 
/* out0282_had-eta2-phi14*/	1, 134, 4, 
/* out0283_had-eta3-phi14*/	2, 133, 3, 134, 2, 
/* out0284_had-eta4-phi14*/	1, 133, 4, 
/* out0285_had-eta5-phi14*/	2, 132, 4, 133, 1, 
/* out0286_had-eta6-phi14*/	1, 132, 4, 
/* out0287_had-eta7-phi14*/	0, 
/* out0288_had-eta8-phi14*/	1, 14, 2, 
/* out0289_had-eta9-phi14*/	4, 14, 7, 70, 3, 74, 1, 75, 7, 
/* out0290_had-eta10-phi14*/	3, 12, 3, 14, 3, 74, 5, 
/* out0291_had-eta11-phi14*/	3, 12, 5, 73, 2, 74, 3, 
/* out0292_had-eta12-phi14*/	4, 10, 1, 12, 1, 17, 2, 73, 4, 
/* out0293_had-eta13-phi14*/	3, 10, 2, 17, 1, 73, 3, 
/* out0294_had-eta14-phi14*/	3, 10, 1, 16, 2, 72, 3, 
/* out0295_had-eta15-phi14*/	2, 16, 2, 72, 2, 
/* out0296_had-eta16-phi14*/	4, 15, 2, 16, 1, 72, 1, 76, 1, 
/* out0297_had-eta17-phi14*/	3, 15, 3, 71, 1, 76, 1, 
/* out0298_had-eta18-phi14*/	2, 15, 1, 71, 1, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	1, 135, 2, 
/* out0301_had-eta1-phi15*/	2, 134, 2, 135, 6, 
/* out0302_had-eta2-phi15*/	1, 134, 4, 
/* out0303_had-eta3-phi15*/	2, 133, 3, 134, 2, 
/* out0304_had-eta4-phi15*/	1, 133, 4, 
/* out0305_had-eta5-phi15*/	2, 132, 4, 133, 1, 
/* out0306_had-eta6-phi15*/	1, 132, 4, 
/* out0307_had-eta7-phi15*/	0, 
/* out0308_had-eta8-phi15*/	0, 
/* out0309_had-eta9-phi15*/	3, 13, 3, 14, 2, 70, 8, 
/* out0310_had-eta10-phi15*/	5, 12, 2, 13, 3, 68, 3, 70, 3, 74, 1, 
/* out0311_had-eta11-phi15*/	2, 12, 4, 68, 4, 
/* out0312_had-eta12-phi15*/	5, 10, 3, 12, 1, 67, 1, 68, 1, 73, 3, 
/* out0313_had-eta13-phi15*/	4, 10, 3, 67, 1, 72, 1, 73, 1, 
/* out0314_had-eta14-phi15*/	3, 9, 1, 10, 2, 72, 3, 
/* out0315_had-eta15-phi15*/	2, 9, 2, 72, 2, 
/* out0316_had-eta16-phi15*/	3, 9, 2, 71, 1, 72, 1, 
/* out0317_had-eta17-phi15*/	2, 15, 3, 71, 2, 
/* out0318_had-eta18-phi15*/	1, 71, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	1, 139, 2, 
/* out0321_had-eta1-phi16*/	2, 138, 2, 139, 6, 
/* out0322_had-eta2-phi16*/	1, 138, 4, 
/* out0323_had-eta3-phi16*/	2, 137, 3, 138, 2, 
/* out0324_had-eta4-phi16*/	1, 137, 4, 
/* out0325_had-eta5-phi16*/	2, 136, 4, 137, 1, 
/* out0326_had-eta6-phi16*/	1, 136, 4, 
/* out0327_had-eta7-phi16*/	0, 
/* out0328_had-eta8-phi16*/	0, 
/* out0329_had-eta9-phi16*/	3, 13, 5, 69, 4, 70, 2, 
/* out0330_had-eta10-phi16*/	4, 11, 1, 13, 5, 68, 3, 69, 3, 
/* out0331_had-eta11-phi16*/	2, 11, 5, 68, 5, 
/* out0332_had-eta12-phi16*/	3, 10, 1, 11, 3, 67, 4, 
/* out0333_had-eta13-phi16*/	3, 10, 2, 48, 1, 67, 3, 
/* out0334_had-eta14-phi16*/	5, 9, 2, 10, 1, 61, 1, 67, 1, 72, 1, 
/* out0335_had-eta15-phi16*/	3, 9, 2, 61, 1, 72, 1, 
/* out0336_had-eta16-phi16*/	2, 9, 2, 71, 2, 
/* out0337_had-eta17-phi16*/	2, 9, 1, 71, 2, 
/* out0338_had-eta18-phi16*/	1, 71, 2, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	1, 139, 2, 
/* out0341_had-eta1-phi17*/	2, 138, 2, 139, 6, 
/* out0342_had-eta2-phi17*/	1, 138, 4, 
/* out0343_had-eta3-phi17*/	2, 137, 3, 138, 2, 
/* out0344_had-eta4-phi17*/	1, 137, 4, 
/* out0345_had-eta5-phi17*/	2, 136, 4, 137, 1, 
/* out0346_had-eta6-phi17*/	1, 136, 4, 
/* out0347_had-eta7-phi17*/	0, 
/* out0348_had-eta8-phi17*/	0, 
/* out0349_had-eta9-phi17*/	2, 51, 3, 69, 5, 
/* out0350_had-eta10-phi17*/	4, 11, 1, 51, 4, 65, 2, 69, 4, 
/* out0351_had-eta11-phi17*/	2, 11, 4, 65, 5, 
/* out0352_had-eta12-phi17*/	4, 11, 2, 48, 1, 65, 1, 67, 3, 
/* out0353_had-eta13-phi17*/	2, 48, 3, 67, 3, 
/* out0354_had-eta14-phi17*/	2, 48, 2, 61, 2, 
/* out0355_had-eta15-phi17*/	2, 9, 2, 61, 2, 
/* out0356_had-eta16-phi17*/	2, 9, 2, 61, 2, 
/* out0357_had-eta17-phi17*/	1, 71, 2, 
/* out0358_had-eta18-phi17*/	1, 71, 2, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	1, 143, 2, 
/* out0361_had-eta1-phi18*/	2, 142, 2, 143, 6, 
/* out0362_had-eta2-phi18*/	1, 142, 4, 
/* out0363_had-eta3-phi18*/	2, 141, 3, 142, 2, 
/* out0364_had-eta4-phi18*/	1, 141, 4, 
/* out0365_had-eta5-phi18*/	2, 140, 4, 141, 1, 
/* out0366_had-eta6-phi18*/	1, 140, 4, 
/* out0367_had-eta7-phi18*/	0, 
/* out0368_had-eta8-phi18*/	0, 
/* out0369_had-eta9-phi18*/	2, 51, 4, 66, 5, 
/* out0370_had-eta10-phi18*/	4, 49, 1, 51, 5, 65, 2, 66, 4, 
/* out0371_had-eta11-phi18*/	2, 49, 4, 65, 5, 
/* out0372_had-eta12-phi18*/	4, 48, 2, 49, 2, 62, 3, 65, 1, 
/* out0373_had-eta13-phi18*/	2, 48, 3, 62, 3, 
/* out0374_had-eta14-phi18*/	2, 48, 2, 61, 2, 
/* out0375_had-eta15-phi18*/	2, 5, 2, 61, 2, 
/* out0376_had-eta16-phi18*/	2, 5, 2, 61, 2, 
/* out0377_had-eta17-phi18*/	1, 56, 2, 
/* out0378_had-eta18-phi18*/	1, 56, 2, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	1, 143, 2, 
/* out0381_had-eta1-phi19*/	2, 142, 2, 143, 6, 
/* out0382_had-eta2-phi19*/	1, 142, 4, 
/* out0383_had-eta3-phi19*/	2, 141, 3, 142, 2, 
/* out0384_had-eta4-phi19*/	1, 141, 4, 
/* out0385_had-eta5-phi19*/	2, 140, 4, 141, 1, 
/* out0386_had-eta6-phi19*/	1, 140, 4, 
/* out0387_had-eta7-phi19*/	0, 
/* out0388_had-eta8-phi19*/	0, 
/* out0389_had-eta9-phi19*/	3, 50, 5, 64, 2, 66, 4, 
/* out0390_had-eta10-phi19*/	4, 49, 1, 50, 5, 63, 3, 66, 3, 
/* out0391_had-eta11-phi19*/	2, 49, 5, 63, 5, 
/* out0392_had-eta12-phi19*/	3, 6, 1, 49, 3, 62, 4, 
/* out0393_had-eta13-phi19*/	3, 6, 2, 48, 1, 62, 3, 
/* out0394_had-eta14-phi19*/	6, 5, 2, 6, 1, 48, 1, 57, 1, 61, 1, 62, 1, 
/* out0395_had-eta15-phi19*/	3, 5, 2, 57, 1, 61, 1, 
/* out0396_had-eta16-phi19*/	2, 5, 2, 56, 2, 
/* out0397_had-eta17-phi19*/	2, 5, 1, 56, 2, 
/* out0398_had-eta18-phi19*/	1, 56, 2, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	1, 147, 2, 
/* out0401_had-eta1-phi20*/	2, 146, 2, 147, 6, 
/* out0402_had-eta2-phi20*/	1, 146, 4, 
/* out0403_had-eta3-phi20*/	2, 145, 3, 146, 2, 
/* out0404_had-eta4-phi20*/	1, 145, 4, 
/* out0405_had-eta5-phi20*/	2, 144, 4, 145, 1, 
/* out0406_had-eta6-phi20*/	1, 144, 4, 
/* out0407_had-eta7-phi20*/	0, 
/* out0408_had-eta8-phi20*/	0, 
/* out0409_had-eta9-phi20*/	3, 8, 2, 50, 3, 64, 8, 
/* out0410_had-eta10-phi20*/	5, 7, 2, 50, 3, 59, 1, 63, 3, 64, 3, 
/* out0411_had-eta11-phi20*/	2, 7, 4, 63, 4, 
/* out0412_had-eta12-phi20*/	5, 6, 3, 7, 1, 58, 3, 62, 1, 63, 1, 
/* out0413_had-eta13-phi20*/	4, 6, 3, 57, 1, 58, 1, 62, 1, 
/* out0414_had-eta14-phi20*/	3, 5, 1, 6, 2, 57, 3, 
/* out0415_had-eta15-phi20*/	2, 5, 2, 57, 2, 
/* out0416_had-eta16-phi20*/	3, 5, 2, 56, 1, 57, 1, 
/* out0417_had-eta17-phi20*/	2, 0, 3, 56, 2, 
/* out0418_had-eta18-phi20*/	1, 56, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	1, 147, 2, 
/* out0421_had-eta1-phi21*/	2, 146, 2, 147, 6, 
/* out0422_had-eta2-phi21*/	1, 146, 4, 
/* out0423_had-eta3-phi21*/	2, 145, 3, 146, 2, 
/* out0424_had-eta4-phi21*/	1, 145, 4, 
/* out0425_had-eta5-phi21*/	2, 144, 4, 145, 1, 
/* out0426_had-eta6-phi21*/	1, 144, 4, 
/* out0427_had-eta7-phi21*/	0, 
/* out0428_had-eta8-phi21*/	1, 8, 2, 
/* out0429_had-eta9-phi21*/	4, 8, 7, 59, 1, 60, 7, 64, 3, 
/* out0430_had-eta10-phi21*/	3, 7, 3, 8, 3, 59, 5, 
/* out0431_had-eta11-phi21*/	3, 7, 5, 58, 2, 59, 3, 
/* out0432_had-eta12-phi21*/	4, 2, 2, 6, 1, 7, 1, 58, 4, 
/* out0433_had-eta13-phi21*/	3, 2, 1, 6, 2, 58, 3, 
/* out0434_had-eta14-phi21*/	3, 1, 2, 6, 1, 57, 3, 
/* out0435_had-eta15-phi21*/	2, 1, 2, 57, 2, 
/* out0436_had-eta16-phi21*/	4, 0, 2, 1, 1, 52, 1, 57, 1, 
/* out0437_had-eta17-phi21*/	3, 0, 3, 52, 1, 56, 1, 
/* out0438_had-eta18-phi21*/	2, 0, 1, 56, 1, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	1, 151, 2, 
/* out0441_had-eta1-phi22*/	2, 150, 2, 151, 6, 
/* out0442_had-eta2-phi22*/	1, 150, 4, 
/* out0443_had-eta3-phi22*/	2, 149, 3, 150, 2, 
/* out0444_had-eta4-phi22*/	1, 149, 4, 
/* out0445_had-eta5-phi22*/	2, 148, 4, 149, 1, 
/* out0446_had-eta6-phi22*/	1, 148, 4, 
/* out0447_had-eta7-phi22*/	0, 
/* out0448_had-eta8-phi22*/	1, 4, 1, 
/* out0449_had-eta9-phi22*/	5, 3, 1, 4, 7, 8, 2, 55, 2, 60, 9, 
/* out0450_had-eta10-phi22*/	3, 3, 5, 55, 2, 59, 4, 
/* out0451_had-eta11-phi22*/	4, 2, 1, 3, 3, 54, 3, 59, 2, 
/* out0452_had-eta12-phi22*/	3, 2, 4, 54, 2, 58, 2, 
/* out0453_had-eta13-phi22*/	3, 2, 3, 53, 3, 58, 1, 
/* out0454_had-eta14-phi22*/	2, 1, 3, 53, 3, 
/* out0455_had-eta15-phi22*/	4, 1, 2, 52, 2, 53, 1, 57, 1, 
/* out0456_had-eta16-phi22*/	3, 0, 1, 1, 1, 52, 2, 
/* out0457_had-eta17-phi22*/	2, 0, 3, 52, 2, 
/* out0458_had-eta18-phi22*/	2, 0, 1, 52, 1, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	1, 151, 2, 
/* out0461_had-eta1-phi23*/	2, 150, 2, 151, 6, 
/* out0462_had-eta2-phi23*/	1, 150, 4, 
/* out0463_had-eta3-phi23*/	2, 149, 3, 150, 2, 
/* out0464_had-eta4-phi23*/	1, 149, 4, 
/* out0465_had-eta5-phi23*/	2, 148, 4, 149, 1, 
/* out0466_had-eta6-phi23*/	1, 148, 4, 
/* out0467_had-eta7-phi23*/	0, 
/* out0468_had-eta8-phi23*/	0, 
/* out0469_had-eta9-phi23*/	3, 3, 1, 4, 8, 55, 6, 
/* out0470_had-eta10-phi23*/	2, 3, 4, 55, 6, 
/* out0471_had-eta11-phi23*/	2, 3, 2, 54, 6, 
/* out0472_had-eta12-phi23*/	2, 2, 3, 54, 5, 
/* out0473_had-eta13-phi23*/	2, 2, 2, 53, 4, 
/* out0474_had-eta14-phi23*/	2, 1, 2, 53, 3, 
/* out0475_had-eta15-phi23*/	3, 1, 2, 52, 2, 53, 2, 
/* out0476_had-eta16-phi23*/	2, 1, 1, 52, 2, 
/* out0477_had-eta17-phi23*/	2, 0, 1, 52, 2, 
/* out0478_had-eta18-phi23*/	2, 0, 1, 52, 1, 
/* out0479_had-eta19-phi23*/	0, 
};