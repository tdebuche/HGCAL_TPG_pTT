parameter integer matrixH [0:6279] = {
/* num inputs = 166(in0-in165) */
/* num outputs = 480(out0-out479 */
//* max inputs per outputs = 10 */
//* total number of input in adders 1933 */

/* out0000_had-eta0-phi0*/	1, 121, 0, 2, 
/* out0001_had-eta1-phi0*/	1, 121, 0, 4, 
/* out0002_had-eta2-phi0*/	2, 120, 0, 3, 121, 0, 2, 
/* out0003_had-eta3-phi0*/	3, 36, 1, 9, 36, 2, 11, 120, 0, 4, 
/* out0004_had-eta4-phi0*/	7, 27, 0, 1, 27, 2, 3, 35, 1, 5, 35, 2, 9, 36, 1, 1, 119, 0, 3, 120, 0, 1, 
/* out0005_had-eta5-phi0*/	6, 27, 0, 15, 27, 1, 15, 27, 2, 13, 34, 2, 6, 35, 1, 3, 119, 0, 4, 
/* out0006_had-eta6-phi0*/	8, 26, 0, 11, 26, 1, 1, 26, 2, 16, 27, 1, 1, 34, 1, 5, 34, 2, 1, 118, 0, 3, 119, 0, 1, 
/* out0007_had-eta7-phi0*/	7, 25, 0, 2, 25, 2, 3, 26, 0, 5, 26, 1, 15, 33, 1, 2, 33, 2, 4, 118, 0, 3, 
/* out0008_had-eta8-phi0*/	5, 25, 0, 12, 25, 1, 2, 25, 2, 13, 33, 1, 1, 118, 0, 2, 
/* out0009_had-eta9-phi0*/	6, 24, 0, 2, 24, 2, 14, 25, 0, 2, 25, 1, 14, 32, 1, 1, 32, 2, 2, 
/* out0010_had-eta10-phi0*/	3, 24, 0, 9, 24, 1, 1, 24, 2, 2, 
/* out0011_had-eta11-phi0*/	7, 3, 3, 2, 3, 8, 16, 3, 9, 7, 9, 5, 2, 9, 11, 2, 24, 0, 3, 24, 1, 15, 
/* out0012_had-eta12-phi0*/	5, 3, 0, 1, 3, 2, 8, 3, 3, 12, 3, 9, 9, 3, 10, 5, 
/* out0013_had-eta13-phi0*/	5, 3, 1, 9, 3, 2, 8, 3, 6, 16, 3, 7, 4, 3, 10, 11, 
/* out0014_had-eta14-phi0*/	6, 1, 3, 2, 1, 8, 16, 1, 9, 9, 3, 1, 2, 3, 4, 16, 3, 7, 12, 
/* out0015_had-eta15-phi0*/	4, 1, 2, 5, 1, 3, 5, 1, 9, 7, 1, 10, 15, 
/* out0016_had-eta16-phi0*/	4, 1, 1, 1, 1, 2, 11, 1, 6, 3, 1, 10, 1, 
/* out0017_had-eta17-phi0*/	3, 1, 1, 2, 1, 6, 13, 1, 7, 9, 
/* out0018_had-eta18-phi0*/	4, 0, 3, 16, 0, 4, 8, 1, 4, 16, 1, 7, 5, 
/* out0019_had-eta19-phi0*/	4, 0, 1, 9, 0, 2, 1, 0, 4, 4, 0, 5, 16, 
/* out0020_had-eta0-phi1*/	1, 121, 0, 2, 
/* out0021_had-eta1-phi1*/	1, 121, 0, 4, 
/* out0022_had-eta2-phi1*/	4, 36, 2, 1, 47, 1, 3, 120, 0, 3, 121, 0, 2, 
/* out0023_had-eta3-phi1*/	6, 36, 0, 16, 36, 1, 5, 36, 2, 4, 46, 2, 9, 47, 1, 9, 120, 0, 4, 
/* out0024_had-eta4-phi1*/	8, 35, 0, 15, 35, 1, 3, 35, 2, 7, 36, 1, 1, 45, 2, 2, 46, 1, 7, 119, 0, 3, 120, 0, 1, 
/* out0025_had-eta5-phi1*/	7, 34, 0, 8, 34, 2, 9, 35, 0, 1, 35, 1, 5, 45, 1, 2, 45, 2, 2, 119, 0, 4, 
/* out0026_had-eta6-phi1*/	6, 33, 0, 1, 33, 2, 5, 34, 0, 6, 34, 1, 11, 118, 0, 3, 119, 0, 1, 
/* out0027_had-eta7-phi1*/	4, 33, 0, 7, 33, 1, 6, 33, 2, 7, 118, 0, 3, 
/* out0028_had-eta8-phi1*/	3, 32, 2, 8, 33, 1, 7, 118, 0, 2, 
/* out0029_had-eta9-phi1*/	3, 32, 0, 1, 32, 1, 8, 32, 2, 5, 
/* out0030_had-eta10-phi1*/	4, 9, 8, 15, 9, 9, 4, 24, 0, 2, 32, 1, 4, 
/* out0031_had-eta11-phi1*/	5, 9, 5, 8, 9, 6, 6, 9, 8, 1, 9, 10, 9, 9, 11, 14, 
/* out0032_had-eta12-phi1*/	6, 3, 0, 8, 3, 3, 2, 8, 8, 1, 9, 4, 12, 9, 5, 6, 9, 6, 1, 
/* out0033_had-eta13-phi1*/	4, 3, 0, 7, 3, 1, 4, 8, 8, 9, 8, 11, 7, 
/* out0034_had-eta14-phi1*/	4, 1, 3, 2, 3, 1, 1, 8, 5, 10, 8, 11, 8, 
/* out0035_had-eta15-phi1*/	4, 1, 0, 6, 1, 3, 7, 8, 4, 3, 8, 5, 3, 
/* out0036_had-eta16-phi1*/	3, 1, 0, 9, 1, 1, 5, 2, 8, 1, 
/* out0037_had-eta17-phi1*/	3, 1, 1, 8, 1, 7, 1, 2, 11, 5, 
/* out0038_had-eta18-phi1*/	5, 0, 2, 4, 0, 4, 4, 1, 7, 1, 2, 5, 3, 2, 11, 1, 
/* out0039_had-eta19-phi1*/	3, 0, 0, 1, 0, 1, 7, 0, 2, 10, 
/* out0040_had-eta0-phi2*/	1, 125, 0, 2, 
/* out0041_had-eta1-phi2*/	1, 125, 0, 4, 
/* out0042_had-eta2-phi2*/	4, 47, 0, 10, 58, 2, 6, 124, 0, 3, 125, 0, 2, 
/* out0043_had-eta3-phi2*/	8, 46, 0, 11, 46, 2, 7, 47, 0, 6, 47, 1, 4, 57, 2, 1, 58, 1, 9, 58, 2, 8, 124, 0, 4, 
/* out0044_had-eta4-phi2*/	8, 45, 0, 6, 45, 2, 9, 46, 0, 5, 46, 1, 9, 57, 1, 2, 57, 2, 4, 123, 0, 3, 124, 0, 1, 
/* out0045_had-eta5-phi2*/	6, 34, 0, 1, 44, 2, 4, 45, 0, 7, 45, 1, 14, 45, 2, 3, 123, 0, 4, 
/* out0046_had-eta6-phi2*/	6, 34, 0, 1, 44, 0, 3, 44, 1, 8, 44, 2, 12, 122, 0, 3, 123, 0, 1, 
/* out0047_had-eta7-phi2*/	4, 33, 0, 7, 43, 2, 8, 44, 1, 5, 122, 0, 3, 
/* out0048_had-eta8-phi2*/	6, 32, 0, 4, 32, 2, 1, 33, 0, 1, 43, 1, 7, 43, 2, 3, 122, 0, 2, 
/* out0049_had-eta9-phi2*/	3, 32, 0, 10, 32, 1, 1, 42, 2, 2, 
/* out0050_had-eta10-phi2*/	8, 9, 2, 1, 9, 3, 13, 9, 9, 12, 9, 10, 2, 32, 0, 1, 32, 1, 2, 42, 1, 1, 42, 2, 1, 
/* out0051_had-eta11-phi2*/	6, 9, 0, 2, 9, 1, 5, 9, 2, 15, 9, 3, 3, 9, 6, 7, 9, 10, 5, 
/* out0052_had-eta12-phi2*/	6, 8, 8, 2, 8, 9, 5, 9, 1, 2, 9, 4, 4, 9, 6, 2, 9, 7, 15, 
/* out0053_had-eta13-phi2*/	5, 8, 2, 1, 8, 8, 4, 8, 9, 9, 8, 10, 11, 8, 11, 1, 
/* out0054_had-eta14-phi2*/	4, 8, 2, 1, 8, 5, 2, 8, 6, 13, 8, 10, 5, 
/* out0055_had-eta15-phi2*/	4, 2, 8, 1, 8, 4, 13, 8, 5, 1, 8, 7, 3, 
/* out0056_had-eta16-phi2*/	3, 1, 0, 1, 2, 8, 13, 2, 11, 1, 
/* out0057_had-eta17-phi2*/	2, 2, 10, 3, 2, 11, 9, 
/* out0058_had-eta18-phi2*/	2, 2, 5, 9, 2, 6, 1, 
/* out0059_had-eta19-phi2*/	4, 0, 0, 15, 0, 2, 1, 2, 4, 4, 2, 5, 2, 
/* out0060_had-eta0-phi3*/	1, 125, 0, 2, 
/* out0061_had-eta1-phi3*/	1, 125, 0, 4, 
/* out0062_had-eta2-phi3*/	5, 58, 0, 2, 58, 2, 1, 100, 2, 1, 124, 0, 3, 125, 0, 2, 
/* out0063_had-eta3-phi3*/	8, 57, 0, 4, 57, 2, 6, 58, 0, 14, 58, 1, 7, 58, 2, 1, 100, 1, 5, 100, 2, 9, 124, 0, 4, 
/* out0064_had-eta4-phi3*/	8, 45, 0, 1, 56, 0, 1, 56, 2, 3, 57, 0, 11, 57, 1, 14, 57, 2, 5, 123, 0, 3, 124, 0, 1, 
/* out0065_had-eta5-phi3*/	6, 44, 0, 1, 45, 0, 2, 56, 0, 2, 56, 1, 10, 56, 2, 13, 123, 0, 4, 
/* out0066_had-eta6-phi3*/	6, 44, 0, 12, 44, 1, 1, 55, 2, 8, 56, 1, 3, 122, 0, 3, 123, 0, 1, 
/* out0067_had-eta7-phi3*/	5, 43, 0, 8, 43, 2, 5, 44, 1, 2, 55, 1, 4, 122, 0, 3, 
/* out0068_had-eta8-phi3*/	4, 42, 2, 1, 43, 0, 6, 43, 1, 9, 122, 0, 2, 
/* out0069_had-eta9-phi3*/	2, 42, 0, 1, 42, 2, 11, 
/* out0070_had-eta10-phi3*/	3, 9, 0, 2, 42, 1, 10, 42, 2, 1, 
/* out0071_had-eta11-phi3*/	5, 9, 0, 12, 9, 1, 4, 10, 8, 13, 10, 11, 5, 42, 1, 1, 
/* out0072_had-eta12-phi3*/	6, 8, 3, 3, 8, 9, 2, 9, 1, 5, 9, 7, 1, 10, 5, 10, 10, 11, 10, 
/* out0073_had-eta13-phi3*/	4, 8, 0, 6, 8, 2, 6, 8, 3, 13, 10, 5, 1, 
/* out0074_had-eta14-phi3*/	5, 8, 0, 1, 8, 1, 9, 8, 2, 8, 8, 6, 3, 8, 7, 1, 
/* out0075_had-eta15-phi3*/	3, 2, 9, 5, 8, 1, 1, 8, 7, 12, 
/* out0076_had-eta16-phi3*/	3, 2, 8, 1, 2, 9, 10, 2, 10, 4, 
/* out0077_had-eta17-phi3*/	3, 2, 2, 1, 2, 6, 3, 2, 10, 9, 
/* out0078_had-eta18-phi3*/	4, 2, 4, 1, 2, 5, 2, 2, 6, 8, 2, 7, 1, 
/* out0079_had-eta19-phi3*/	2, 2, 4, 9, 2, 7, 1, 
/* out0080_had-eta0-phi4*/	1, 129, 0, 2, 
/* out0081_had-eta1-phi4*/	1, 129, 0, 4, 
/* out0082_had-eta2-phi4*/	4, 100, 0, 2, 100, 2, 2, 128, 0, 3, 129, 0, 2, 
/* out0083_had-eta3-phi4*/	8, 99, 0, 1, 99, 2, 2, 100, 0, 14, 100, 1, 11, 100, 2, 4, 101, 1, 1, 101, 2, 5, 128, 0, 4, 
/* out0084_had-eta4-phi4*/	7, 56, 0, 1, 57, 0, 1, 99, 0, 7, 99, 1, 12, 99, 2, 14, 127, 0, 3, 128, 0, 1, 
/* out0085_had-eta5-phi4*/	6, 56, 0, 12, 56, 1, 2, 98, 1, 2, 98, 2, 10, 99, 1, 2, 127, 0, 4, 
/* out0086_had-eta6-phi4*/	7, 55, 0, 11, 55, 1, 1, 55, 2, 8, 56, 1, 1, 98, 1, 2, 126, 0, 3, 127, 0, 1, 
/* out0087_had-eta7-phi4*/	5, 43, 0, 1, 54, 2, 6, 55, 0, 2, 55, 1, 11, 126, 0, 3, 
/* out0088_had-eta8-phi4*/	5, 42, 0, 1, 43, 0, 1, 54, 1, 6, 54, 2, 9, 126, 0, 2, 
/* out0089_had-eta9-phi4*/	2, 42, 0, 10, 54, 1, 2, 
/* out0090_had-eta10-phi4*/	5, 10, 3, 2, 10, 9, 4, 42, 0, 4, 42, 1, 4, 64, 2, 1, 
/* out0091_had-eta11-phi4*/	6, 10, 2, 6, 10, 3, 4, 10, 8, 3, 10, 9, 12, 10, 10, 12, 10, 11, 1, 
/* out0092_had-eta12-phi4*/	6, 10, 2, 2, 10, 4, 2, 10, 5, 5, 10, 6, 15, 10, 7, 3, 10, 10, 4, 
/* out0093_had-eta13-phi4*/	3, 8, 0, 6, 10, 4, 13, 14, 8, 5, 
/* out0094_had-eta14-phi4*/	4, 8, 0, 3, 8, 1, 4, 14, 8, 5, 14, 11, 7, 
/* out0095_had-eta15-phi4*/	5, 2, 3, 4, 2, 9, 1, 8, 1, 2, 14, 5, 6, 14, 11, 4, 
/* out0096_had-eta16-phi4*/	2, 2, 2, 2, 2, 3, 12, 
/* out0097_had-eta17-phi4*/	2, 2, 1, 1, 2, 2, 11, 
/* out0098_had-eta18-phi4*/	4, 2, 1, 1, 2, 2, 2, 2, 6, 4, 2, 7, 4, 
/* out0099_had-eta19-phi4*/	2, 2, 4, 2, 2, 7, 6, 
/* out0100_had-eta0-phi5*/	1, 129, 0, 2, 
/* out0101_had-eta1-phi5*/	1, 129, 0, 4, 
/* out0102_had-eta2-phi5*/	3, 101, 2, 1, 128, 0, 3, 129, 0, 2, 
/* out0103_had-eta3-phi5*/	5, 101, 0, 16, 101, 1, 13, 101, 2, 10, 108, 2, 1, 128, 0, 4, 
/* out0104_had-eta4-phi5*/	7, 99, 0, 8, 99, 1, 2, 101, 1, 2, 108, 1, 6, 108, 2, 15, 127, 0, 3, 128, 0, 1, 
/* out0105_had-eta5-phi5*/	5, 98, 0, 16, 98, 1, 5, 98, 2, 6, 108, 1, 2, 127, 0, 4, 
/* out0106_had-eta6-phi5*/	5, 55, 0, 2, 98, 1, 7, 106, 2, 13, 126, 0, 3, 127, 0, 1, 
/* out0107_had-eta7-phi5*/	6, 54, 0, 6, 54, 2, 1, 55, 0, 1, 106, 1, 8, 106, 2, 3, 126, 0, 3, 
/* out0108_had-eta8-phi5*/	3, 54, 0, 10, 54, 1, 5, 126, 0, 2, 
/* out0109_had-eta9-phi5*/	2, 54, 1, 3, 64, 2, 10, 
/* out0110_had-eta10-phi5*/	3, 10, 3, 1, 64, 1, 6, 64, 2, 5, 
/* out0111_had-eta11-phi5*/	5, 10, 0, 15, 10, 1, 2, 10, 2, 4, 10, 3, 9, 64, 1, 1, 
/* out0112_had-eta12-phi5*/	5, 10, 0, 1, 10, 1, 14, 10, 2, 4, 10, 6, 1, 10, 7, 9, 
/* out0113_had-eta13-phi5*/	5, 10, 4, 1, 10, 7, 4, 14, 8, 5, 14, 9, 15, 14, 10, 1, 
/* out0114_had-eta14-phi5*/	4, 14, 6, 2, 14, 8, 1, 14, 10, 14, 14, 11, 4, 
/* out0115_had-eta15-phi5*/	4, 14, 4, 2, 14, 5, 10, 14, 6, 5, 14, 11, 1, 
/* out0116_had-eta16-phi5*/	2, 2, 0, 9, 14, 4, 5, 
/* out0117_had-eta17-phi5*/	2, 2, 0, 7, 2, 1, 5, 
/* out0118_had-eta18-phi5*/	2, 2, 1, 9, 2, 7, 1, 
/* out0119_had-eta19-phi5*/	1, 2, 7, 3, 
/* out0120_had-eta0-phi6*/	1, 133, 0, 2, 
/* out0121_had-eta1-phi6*/	1, 133, 0, 4, 
/* out0122_had-eta2-phi6*/	3, 110, 0, 1, 132, 0, 3, 133, 0, 2, 
/* out0123_had-eta3-phi6*/	5, 108, 0, 1, 110, 0, 10, 110, 1, 13, 110, 2, 16, 132, 0, 4, 
/* out0124_had-eta4-phi6*/	7, 108, 0, 15, 108, 1, 6, 109, 1, 2, 109, 2, 8, 110, 1, 2, 131, 0, 3, 132, 0, 1, 
/* out0125_had-eta5-phi6*/	5, 107, 0, 6, 107, 1, 5, 107, 2, 16, 108, 1, 2, 131, 0, 4, 
/* out0126_had-eta6-phi6*/	5, 66, 2, 2, 106, 0, 13, 107, 1, 7, 130, 0, 3, 131, 0, 1, 
/* out0127_had-eta7-phi6*/	6, 65, 0, 1, 65, 2, 6, 66, 2, 1, 106, 0, 3, 106, 1, 8, 130, 0, 3, 
/* out0128_had-eta8-phi6*/	3, 65, 1, 5, 65, 2, 10, 130, 0, 2, 
/* out0129_had-eta9-phi6*/	2, 64, 0, 10, 65, 1, 3, 
/* out0130_had-eta10-phi6*/	3, 15, 9, 1, 64, 0, 4, 64, 1, 7, 
/* out0131_had-eta11-phi6*/	5, 15, 8, 15, 15, 9, 9, 15, 10, 4, 15, 11, 2, 64, 1, 2, 
/* out0132_had-eta12-phi6*/	5, 15, 5, 9, 15, 6, 1, 15, 8, 1, 15, 10, 4, 15, 11, 14, 
/* out0133_had-eta13-phi6*/	6, 14, 0, 3, 14, 2, 2, 14, 3, 15, 14, 9, 1, 15, 4, 1, 15, 5, 4, 
/* out0134_had-eta14-phi6*/	6, 14, 0, 1, 14, 1, 3, 14, 2, 14, 14, 3, 1, 14, 6, 3, 14, 10, 1, 
/* out0135_had-eta15-phi6*/	3, 14, 4, 3, 14, 6, 6, 14, 7, 9, 
/* out0136_had-eta16-phi6*/	2, 14, 4, 6, 18, 8, 9, 
/* out0137_had-eta17-phi6*/	2, 18, 8, 7, 18, 11, 5, 
/* out0138_had-eta18-phi6*/	2, 18, 5, 1, 18, 11, 9, 
/* out0139_had-eta19-phi6*/	1, 18, 5, 3, 
/* out0140_had-eta0-phi7*/	1, 133, 0, 2, 
/* out0141_had-eta1-phi7*/	1, 133, 0, 4, 
/* out0142_had-eta2-phi7*/	4, 111, 0, 2, 111, 2, 2, 132, 0, 3, 133, 0, 2, 
/* out0143_had-eta3-phi7*/	8, 109, 0, 2, 109, 2, 1, 110, 0, 5, 110, 1, 1, 111, 0, 4, 111, 1, 11, 111, 2, 14, 132, 0, 4, 
/* out0144_had-eta4-phi7*/	7, 67, 2, 1, 68, 2, 1, 109, 0, 14, 109, 1, 12, 109, 2, 7, 131, 0, 3, 132, 0, 1, 
/* out0145_had-eta5-phi7*/	6, 67, 1, 2, 67, 2, 12, 107, 0, 10, 107, 1, 2, 109, 1, 2, 131, 0, 4, 
/* out0146_had-eta6-phi7*/	7, 66, 0, 8, 66, 1, 1, 66, 2, 11, 67, 1, 1, 107, 1, 2, 130, 0, 3, 131, 0, 1, 
/* out0147_had-eta7-phi7*/	5, 65, 0, 6, 66, 1, 11, 66, 2, 2, 77, 2, 1, 130, 0, 3, 
/* out0148_had-eta8-phi7*/	5, 65, 0, 9, 65, 1, 6, 76, 2, 1, 77, 2, 1, 130, 0, 2, 
/* out0149_had-eta9-phi7*/	3, 64, 0, 1, 65, 1, 2, 76, 2, 10, 
/* out0150_had-eta10-phi7*/	5, 15, 3, 4, 15, 9, 2, 64, 0, 1, 76, 1, 4, 76, 2, 4, 
/* out0151_had-eta11-phi7*/	6, 15, 0, 3, 15, 1, 1, 15, 2, 12, 15, 3, 12, 15, 9, 4, 15, 10, 6, 
/* out0152_had-eta12-phi7*/	6, 15, 2, 4, 15, 4, 2, 15, 5, 3, 15, 6, 15, 15, 7, 5, 15, 10, 2, 
/* out0153_had-eta13-phi7*/	3, 14, 0, 7, 15, 4, 13, 19, 8, 6, 
/* out0154_had-eta14-phi7*/	4, 14, 0, 5, 14, 1, 9, 19, 8, 3, 19, 11, 4, 
/* out0155_had-eta15-phi7*/	6, 14, 1, 4, 14, 7, 7, 18, 3, 1, 18, 9, 4, 19, 5, 1, 19, 11, 2, 
/* out0156_had-eta16-phi7*/	2, 18, 9, 12, 18, 10, 2, 
/* out0157_had-eta17-phi7*/	2, 18, 10, 11, 18, 11, 1, 
/* out0158_had-eta18-phi7*/	4, 18, 5, 4, 18, 6, 4, 18, 10, 2, 18, 11, 1, 
/* out0159_had-eta19-phi7*/	2, 18, 4, 2, 18, 5, 6, 
/* out0160_had-eta0-phi8*/	1, 137, 0, 2, 
/* out0161_had-eta1-phi8*/	1, 137, 0, 4, 
/* out0162_had-eta2-phi8*/	5, 69, 0, 1, 69, 2, 2, 111, 0, 1, 136, 0, 3, 137, 0, 2, 
/* out0163_had-eta3-phi8*/	8, 68, 0, 6, 68, 2, 4, 69, 0, 1, 69, 1, 7, 69, 2, 14, 111, 0, 9, 111, 1, 5, 136, 0, 4, 
/* out0164_had-eta4-phi8*/	8, 67, 0, 3, 67, 2, 1, 68, 0, 5, 68, 1, 14, 68, 2, 11, 79, 2, 1, 135, 0, 3, 136, 0, 1, 
/* out0165_had-eta5-phi8*/	6, 67, 0, 13, 67, 1, 10, 67, 2, 2, 78, 2, 1, 79, 2, 2, 135, 0, 4, 
/* out0166_had-eta6-phi8*/	6, 66, 0, 8, 67, 1, 3, 78, 1, 1, 78, 2, 12, 134, 0, 3, 135, 0, 1, 
/* out0167_had-eta7-phi8*/	5, 66, 1, 4, 77, 0, 5, 77, 2, 8, 78, 1, 2, 134, 0, 3, 
/* out0168_had-eta8-phi8*/	4, 76, 0, 1, 77, 1, 9, 77, 2, 6, 134, 0, 2, 
/* out0169_had-eta9-phi8*/	2, 76, 0, 11, 76, 2, 1, 
/* out0170_had-eta10-phi8*/	3, 20, 8, 2, 76, 0, 1, 76, 1, 10, 
/* out0171_had-eta11-phi8*/	5, 15, 0, 13, 15, 1, 5, 20, 8, 13, 20, 11, 4, 76, 1, 1, 
/* out0172_had-eta12-phi8*/	6, 15, 1, 10, 15, 7, 10, 19, 3, 2, 19, 9, 3, 20, 5, 1, 20, 11, 5, 
/* out0173_had-eta13-phi8*/	4, 15, 7, 1, 19, 8, 6, 19, 9, 13, 19, 10, 6, 
/* out0174_had-eta14-phi8*/	5, 19, 5, 1, 19, 6, 3, 19, 8, 1, 19, 10, 8, 19, 11, 9, 
/* out0175_had-eta15-phi8*/	3, 18, 3, 5, 19, 5, 11, 19, 11, 1, 
/* out0176_had-eta16-phi8*/	3, 18, 0, 1, 18, 2, 4, 18, 3, 10, 
/* out0177_had-eta17-phi8*/	3, 18, 2, 9, 18, 6, 3, 18, 10, 1, 
/* out0178_had-eta18-phi8*/	4, 18, 4, 1, 18, 5, 1, 18, 6, 8, 18, 7, 2, 
/* out0179_had-eta19-phi8*/	2, 18, 4, 9, 18, 5, 1, 
/* out0180_had-eta0-phi9*/	1, 137, 0, 2, 
/* out0181_had-eta1-phi9*/	1, 137, 0, 4, 
/* out0182_had-eta2-phi9*/	4, 69, 0, 6, 81, 1, 10, 136, 0, 3, 137, 0, 2, 
/* out0183_had-eta3-phi9*/	8, 68, 0, 1, 69, 0, 8, 69, 1, 9, 80, 0, 7, 80, 2, 11, 81, 0, 4, 81, 1, 6, 136, 0, 4, 
/* out0184_had-eta4-phi9*/	8, 68, 0, 4, 68, 1, 2, 79, 0, 9, 79, 2, 6, 80, 1, 9, 80, 2, 5, 135, 0, 3, 136, 0, 1, 
/* out0185_had-eta5-phi9*/	6, 78, 0, 4, 79, 0, 3, 79, 1, 14, 79, 2, 7, 90, 2, 1, 135, 0, 4, 
/* out0186_had-eta6-phi9*/	6, 78, 0, 12, 78, 1, 8, 78, 2, 3, 90, 2, 1, 134, 0, 3, 135, 0, 1, 
/* out0187_had-eta7-phi9*/	4, 77, 0, 8, 78, 1, 5, 89, 2, 7, 134, 0, 3, 
/* out0188_had-eta8-phi9*/	6, 77, 0, 3, 77, 1, 7, 88, 0, 1, 88, 2, 4, 89, 2, 1, 134, 0, 2, 
/* out0189_had-eta9-phi9*/	3, 76, 0, 2, 88, 1, 1, 88, 2, 10, 
/* out0190_had-eta10-phi9*/	8, 20, 2, 2, 20, 3, 12, 20, 9, 13, 20, 10, 1, 76, 0, 1, 76, 1, 1, 88, 1, 2, 88, 2, 1, 
/* out0191_had-eta11-phi9*/	6, 20, 2, 5, 20, 6, 7, 20, 8, 1, 20, 9, 3, 20, 10, 15, 20, 11, 5, 
/* out0192_had-eta12-phi9*/	6, 19, 0, 2, 19, 3, 5, 20, 4, 4, 20, 5, 15, 20, 6, 2, 20, 11, 2, 
/* out0193_had-eta13-phi9*/	5, 19, 0, 4, 19, 1, 1, 19, 2, 11, 19, 3, 9, 19, 10, 1, 
/* out0194_had-eta14-phi9*/	4, 19, 2, 5, 19, 6, 13, 19, 7, 2, 19, 10, 1, 
/* out0195_had-eta15-phi9*/	4, 18, 0, 1, 19, 4, 13, 19, 5, 3, 19, 7, 1, 
/* out0196_had-eta16-phi9*/	2, 18, 0, 13, 18, 1, 1, 
/* out0197_had-eta17-phi9*/	2, 18, 1, 9, 18, 2, 3, 
/* out0198_had-eta18-phi9*/	2, 18, 6, 1, 18, 7, 9, 
/* out0199_had-eta19-phi9*/	3, 4, 4, 14, 18, 4, 4, 18, 7, 2, 
/* out0200_had-eta0-phi10*/	1, 141, 0, 2, 
/* out0201_had-eta1-phi10*/	1, 141, 0, 4, 
/* out0202_had-eta2-phi10*/	4, 81, 0, 3, 92, 0, 1, 140, 0, 3, 141, 0, 2, 
/* out0203_had-eta3-phi10*/	6, 80, 0, 9, 81, 0, 9, 92, 0, 4, 92, 1, 5, 92, 2, 16, 140, 0, 4, 
/* out0204_had-eta4-phi10*/	8, 79, 0, 2, 80, 1, 7, 91, 0, 7, 91, 1, 3, 91, 2, 15, 92, 1, 1, 139, 0, 3, 140, 0, 1, 
/* out0205_had-eta5-phi10*/	7, 79, 0, 2, 79, 1, 2, 90, 0, 9, 90, 2, 8, 91, 1, 5, 91, 2, 1, 139, 0, 4, 
/* out0206_had-eta6-phi10*/	6, 89, 0, 5, 89, 2, 1, 90, 1, 11, 90, 2, 6, 138, 0, 3, 139, 0, 1, 
/* out0207_had-eta7-phi10*/	4, 89, 0, 7, 89, 1, 6, 89, 2, 7, 138, 0, 3, 
/* out0208_had-eta8-phi10*/	3, 88, 0, 8, 89, 1, 7, 138, 0, 2, 
/* out0209_had-eta9-phi10*/	3, 88, 0, 5, 88, 1, 8, 88, 2, 1, 
/* out0210_had-eta10-phi10*/	4, 20, 0, 15, 20, 3, 4, 28, 2, 1, 88, 1, 4, 
/* out0211_had-eta11-phi10*/	5, 20, 0, 1, 20, 1, 14, 20, 2, 9, 20, 6, 6, 20, 7, 8, 
/* out0212_had-eta12-phi10*/	6, 7, 8, 8, 7, 9, 1, 19, 0, 1, 20, 4, 12, 20, 6, 1, 20, 7, 6, 
/* out0213_had-eta13-phi10*/	4, 7, 8, 6, 7, 11, 3, 19, 0, 9, 19, 1, 7, 
/* out0214_had-eta14-phi10*/	3, 6, 9, 1, 19, 1, 8, 19, 7, 10, 
/* out0215_had-eta15-phi10*/	4, 6, 8, 6, 6, 9, 6, 19, 4, 3, 19, 7, 3, 
/* out0216_had-eta16-phi10*/	3, 6, 8, 10, 6, 11, 4, 18, 0, 1, 
/* out0217_had-eta17-phi10*/	2, 6, 11, 7, 18, 1, 5, 
/* out0218_had-eta18-phi10*/	5, 4, 3, 1, 4, 5, 4, 6, 5, 1, 18, 1, 1, 18, 7, 3, 
/* out0219_had-eta19-phi10*/	3, 4, 4, 2, 4, 5, 10, 4, 6, 6, 
/* out0220_had-eta0-phi11*/	1, 141, 0, 2, 
/* out0221_had-eta1-phi11*/	1, 141, 0, 4, 
/* out0222_had-eta2-phi11*/	2, 140, 0, 3, 141, 0, 2, 
/* out0223_had-eta3-phi11*/	3, 92, 0, 11, 92, 1, 9, 140, 0, 4, 
/* out0224_had-eta4-phi11*/	7, 31, 0, 3, 31, 2, 1, 91, 0, 9, 91, 1, 5, 92, 1, 1, 139, 0, 3, 140, 0, 1, 
/* out0225_had-eta5-phi11*/	6, 31, 0, 1, 31, 1, 3, 31, 2, 15, 90, 0, 6, 91, 1, 3, 139, 0, 4, 
/* out0226_had-eta6-phi11*/	7, 30, 0, 4, 30, 2, 11, 31, 1, 1, 90, 0, 1, 90, 1, 5, 138, 0, 3, 139, 0, 1, 
/* out0227_had-eta7-phi11*/	7, 29, 0, 3, 29, 2, 1, 30, 1, 4, 30, 2, 5, 89, 0, 4, 89, 1, 2, 138, 0, 3, 
/* out0228_had-eta8-phi11*/	5, 29, 0, 1, 29, 1, 1, 29, 2, 13, 89, 1, 1, 138, 0, 2, 
/* out0229_had-eta9-phi11*/	6, 28, 0, 3, 28, 2, 2, 29, 1, 3, 29, 2, 2, 88, 0, 2, 88, 1, 1, 
/* out0230_had-eta10-phi11*/	3, 28, 0, 1, 28, 1, 1, 28, 2, 10, 
/* out0231_had-eta11-phi11*/	6, 7, 3, 6, 7, 9, 2, 20, 1, 2, 20, 7, 2, 28, 1, 3, 28, 2, 3, 
/* out0232_had-eta12-phi11*/	5, 7, 2, 4, 7, 3, 5, 7, 8, 1, 7, 9, 13, 7, 10, 8, 
/* out0233_had-eta13-phi11*/	5, 7, 5, 3, 7, 6, 4, 7, 8, 1, 7, 10, 8, 7, 11, 10, 
/* out0234_had-eta14-phi11*/	4, 6, 3, 8, 6, 9, 2, 7, 5, 9, 7, 11, 3, 
/* out0235_had-eta15-phi11*/	4, 6, 2, 3, 6, 3, 4, 6, 9, 7, 6, 10, 5, 
/* out0236_had-eta16-phi11*/	3, 6, 6, 2, 6, 10, 11, 6, 11, 2, 
/* out0237_had-eta17-phi11*/	3, 6, 5, 8, 6, 6, 2, 6, 11, 3, 
/* out0238_had-eta18-phi11*/	2, 4, 3, 7, 6, 5, 3, 
/* out0239_had-eta19-phi11*/	4, 4, 2, 5, 4, 3, 3, 4, 5, 2, 4, 6, 10, 
/* out0240_had-eta0-phi12*/	1, 145, 0, 2, 
/* out0241_had-eta1-phi12*/	1, 145, 0, 4, 
/* out0242_had-eta2-phi12*/	2, 144, 0, 3, 145, 0, 2, 
/* out0243_had-eta3-phi12*/	4, 41, 0, 3, 41, 1, 2, 41, 2, 16, 144, 0, 4, 
/* out0244_had-eta4-phi12*/	6, 31, 0, 4, 40, 0, 2, 40, 2, 12, 41, 1, 1, 143, 0, 3, 144, 0, 1, 
/* out0245_had-eta5-phi12*/	7, 31, 0, 8, 31, 1, 11, 39, 0, 1, 39, 2, 5, 40, 1, 1, 40, 2, 2, 143, 0, 4, 
/* out0246_had-eta6-phi12*/	6, 30, 0, 12, 30, 1, 3, 31, 1, 1, 39, 2, 6, 142, 0, 3, 143, 0, 1, 
/* out0247_had-eta7-phi12*/	4, 29, 0, 4, 30, 1, 9, 38, 2, 6, 142, 0, 3, 
/* out0248_had-eta8-phi12*/	4, 29, 0, 8, 29, 1, 7, 38, 2, 1, 142, 0, 2, 
/* out0249_had-eta9-phi12*/	3, 28, 0, 5, 29, 1, 5, 37, 2, 3, 
/* out0250_had-eta10-phi12*/	2, 28, 0, 6, 28, 1, 5, 
/* out0251_had-eta11-phi12*/	4, 7, 0, 8, 7, 3, 1, 13, 8, 4, 28, 1, 6, 
/* out0252_had-eta12-phi12*/	4, 7, 0, 7, 7, 1, 8, 7, 2, 12, 7, 3, 4, 
/* out0253_had-eta13-phi12*/	4, 7, 4, 4, 7, 5, 2, 7, 6, 12, 7, 7, 6, 
/* out0254_had-eta14-phi12*/	4, 6, 0, 8, 6, 3, 1, 7, 4, 9, 7, 5, 2, 
/* out0255_had-eta15-phi12*/	4, 6, 0, 4, 6, 1, 3, 6, 2, 9, 6, 3, 3, 
/* out0256_had-eta16-phi12*/	3, 6, 2, 4, 6, 6, 10, 6, 7, 1, 
/* out0257_had-eta17-phi12*/	4, 6, 4, 6, 6, 5, 4, 6, 6, 2, 6, 7, 1, 
/* out0258_had-eta18-phi12*/	3, 4, 0, 6, 4, 3, 2, 6, 4, 3, 
/* out0259_had-eta19-phi12*/	4, 4, 0, 2, 4, 1, 1, 4, 2, 8, 4, 3, 3, 
/* out0260_had-eta0-phi13*/	1, 145, 0, 2, 
/* out0261_had-eta1-phi13*/	1, 145, 0, 4, 
/* out0262_had-eta2-phi13*/	5, 41, 0, 1, 53, 0, 1, 53, 1, 5, 144, 0, 3, 145, 0, 2, 
/* out0263_had-eta3-phi13*/	7, 41, 0, 12, 41, 1, 12, 52, 0, 2, 52, 2, 7, 53, 0, 3, 53, 1, 11, 144, 0, 4, 
/* out0264_had-eta4-phi13*/	8, 40, 0, 14, 40, 1, 9, 40, 2, 2, 41, 1, 1, 51, 2, 2, 52, 2, 7, 143, 0, 3, 144, 0, 1, 
/* out0265_had-eta5-phi13*/	6, 39, 0, 15, 39, 1, 1, 39, 2, 2, 40, 1, 6, 51, 2, 4, 143, 0, 4, 
/* out0266_had-eta6-phi13*/	6, 38, 0, 6, 39, 1, 14, 39, 2, 3, 50, 2, 1, 142, 0, 3, 143, 0, 1, 
/* out0267_had-eta7-phi13*/	4, 38, 0, 7, 38, 1, 5, 38, 2, 7, 142, 0, 3, 
/* out0268_had-eta8-phi13*/	5, 37, 0, 6, 37, 2, 2, 38, 1, 6, 38, 2, 2, 142, 0, 2, 
/* out0269_had-eta9-phi13*/	3, 37, 0, 2, 37, 1, 3, 37, 2, 9, 
/* out0270_had-eta10-phi13*/	6, 13, 3, 12, 13, 9, 7, 28, 0, 1, 28, 1, 1, 37, 1, 3, 37, 2, 2, 
/* out0271_had-eta11-phi13*/	5, 13, 2, 2, 13, 8, 10, 13, 9, 9, 13, 10, 13, 13, 11, 3, 
/* out0272_had-eta12-phi13*/	8, 7, 0, 1, 7, 1, 8, 7, 7, 1, 11, 3, 1, 13, 5, 4, 13, 8, 2, 13, 10, 1, 13, 11, 13, 
/* out0273_had-eta13-phi13*/	5, 7, 4, 2, 7, 7, 9, 11, 3, 1, 11, 8, 1, 11, 9, 12, 
/* out0274_had-eta14-phi13*/	6, 6, 0, 2, 7, 4, 1, 11, 8, 14, 11, 9, 2, 11, 10, 1, 11, 11, 3, 
/* out0275_had-eta15-phi13*/	4, 6, 0, 2, 6, 1, 11, 11, 8, 1, 11, 11, 5, 
/* out0276_had-eta16-phi13*/	2, 6, 1, 2, 6, 7, 12, 
/* out0277_had-eta17-phi13*/	4, 5, 8, 4, 5, 9, 1, 6, 4, 6, 6, 7, 1, 
/* out0278_had-eta18-phi13*/	3, 4, 0, 5, 5, 8, 5, 6, 4, 1, 
/* out0279_had-eta19-phi13*/	3, 4, 0, 3, 4, 1, 10, 4, 2, 3, 
/* out0280_had-eta0-phi14*/	1, 149, 0, 2, 
/* out0281_had-eta1-phi14*/	1, 149, 0, 4, 
/* out0282_had-eta2-phi14*/	5, 53, 0, 5, 63, 0, 4, 63, 2, 2, 148, 0, 3, 149, 0, 2, 
/* out0283_had-eta3-phi14*/	10, 52, 0, 14, 52, 1, 4, 52, 2, 1, 53, 0, 7, 62, 0, 1, 62, 2, 1, 63, 0, 1, 63, 1, 1, 63, 2, 14, 148, 0, 4, 
/* out0284_had-eta4-phi14*/	7, 51, 0, 13, 51, 2, 2, 52, 1, 12, 52, 2, 1, 62, 2, 6, 147, 0, 3, 148, 0, 1, 
/* out0285_had-eta5-phi14*/	5, 50, 0, 4, 51, 0, 2, 51, 1, 14, 51, 2, 8, 147, 0, 4, 
/* out0286_had-eta6-phi14*/	6, 39, 1, 1, 50, 0, 6, 50, 1, 3, 50, 2, 13, 146, 0, 3, 147, 0, 1, 
/* out0287_had-eta7-phi14*/	7, 38, 0, 3, 38, 1, 4, 49, 0, 3, 49, 2, 4, 50, 1, 3, 50, 2, 2, 146, 0, 3, 
/* out0288_had-eta8-phi14*/	4, 37, 0, 5, 38, 1, 1, 49, 2, 10, 146, 0, 2, 
/* out0289_had-eta9-phi14*/	3, 37, 0, 3, 37, 1, 8, 48, 2, 2, 
/* out0290_had-eta10-phi14*/	6, 13, 0, 16, 13, 1, 5, 13, 2, 2, 13, 3, 4, 37, 1, 2, 48, 2, 2, 
/* out0291_had-eta11-phi14*/	5, 13, 1, 4, 13, 2, 12, 13, 6, 13, 13, 7, 5, 13, 10, 2, 
/* out0292_had-eta12-phi14*/	5, 11, 0, 4, 11, 3, 3, 13, 4, 9, 13, 5, 12, 13, 6, 3, 
/* out0293_had-eta13-phi14*/	5, 11, 0, 2, 11, 2, 9, 11, 3, 11, 11, 9, 2, 11, 10, 3, 
/* out0294_had-eta14-phi14*/	4, 11, 2, 1, 11, 6, 6, 11, 10, 12, 11, 11, 2, 
/* out0295_had-eta15-phi14*/	3, 5, 3, 1, 11, 5, 10, 11, 11, 6, 
/* out0296_had-eta16-phi14*/	3, 5, 3, 6, 5, 9, 8, 6, 7, 1, 
/* out0297_had-eta17-phi14*/	3, 5, 8, 2, 5, 9, 7, 5, 10, 3, 
/* out0298_had-eta18-phi14*/	3, 5, 8, 5, 5, 10, 1, 5, 11, 5, 
/* out0299_had-eta19-phi14*/	2, 4, 1, 5, 5, 11, 5, 
/* out0300_had-eta0-phi15*/	1, 149, 0, 2, 
/* out0301_had-eta1-phi15*/	1, 149, 0, 4, 
/* out0302_had-eta2-phi15*/	4, 63, 0, 5, 105, 0, 1, 148, 0, 3, 149, 0, 2, 
/* out0303_had-eta3-phi15*/	6, 62, 0, 10, 63, 0, 6, 63, 1, 15, 105, 0, 2, 105, 2, 12, 148, 0, 4, 
/* out0304_had-eta4-phi15*/	7, 51, 0, 1, 61, 0, 4, 62, 0, 5, 62, 1, 15, 62, 2, 9, 147, 0, 3, 148, 0, 1, 
/* out0305_had-eta5-phi15*/	6, 50, 0, 1, 51, 1, 2, 61, 0, 6, 61, 1, 3, 61, 2, 15, 147, 0, 4, 
/* out0306_had-eta6-phi15*/	8, 50, 0, 5, 50, 1, 8, 60, 0, 2, 60, 2, 6, 61, 1, 2, 61, 2, 1, 146, 0, 3, 147, 0, 1, 
/* out0307_had-eta7-phi15*/	5, 49, 0, 12, 49, 1, 1, 50, 1, 2, 60, 2, 4, 146, 0, 3, 
/* out0308_had-eta8-phi15*/	4, 48, 0, 1, 49, 1, 13, 49, 2, 2, 146, 0, 2, 
/* out0309_had-eta9-phi15*/	2, 48, 0, 8, 48, 2, 5, 
/* out0310_had-eta10-phi15*/	3, 13, 1, 2, 48, 1, 4, 48, 2, 7, 
/* out0311_had-eta11-phi15*/	6, 12, 3, 5, 12, 8, 1, 12, 9, 13, 13, 1, 5, 13, 4, 1, 13, 7, 11, 
/* out0312_had-eta12-phi15*/	5, 11, 0, 5, 12, 8, 15, 12, 9, 2, 12, 11, 2, 13, 4, 6, 
/* out0313_had-eta13-phi15*/	5, 11, 0, 5, 11, 1, 13, 11, 2, 5, 11, 7, 1, 12, 11, 1, 
/* out0314_had-eta14-phi15*/	5, 11, 2, 1, 11, 4, 3, 11, 5, 1, 11, 6, 10, 11, 7, 7, 
/* out0315_had-eta15-phi15*/	4, 5, 0, 4, 5, 3, 1, 11, 4, 8, 11, 5, 5, 
/* out0316_had-eta16-phi15*/	3, 5, 0, 2, 5, 2, 5, 5, 3, 8, 
/* out0317_had-eta17-phi15*/	3, 5, 2, 5, 5, 6, 1, 5, 10, 7, 
/* out0318_had-eta18-phi15*/	4, 5, 5, 1, 5, 6, 3, 5, 10, 5, 5, 11, 2, 
/* out0319_had-eta19-phi15*/	2, 5, 5, 6, 5, 11, 4, 
/* out0320_had-eta0-phi16*/	1, 153, 0, 2, 
/* out0321_had-eta1-phi16*/	1, 153, 0, 4, 
/* out0322_had-eta2-phi16*/	3, 105, 0, 3, 152, 0, 3, 153, 0, 2, 
/* out0323_had-eta3-phi16*/	7, 103, 0, 4, 104, 0, 1, 104, 2, 6, 105, 0, 10, 105, 1, 16, 105, 2, 4, 152, 0, 4, 
/* out0324_had-eta4-phi16*/	7, 61, 0, 1, 62, 1, 1, 103, 0, 10, 103, 1, 7, 103, 2, 15, 151, 0, 3, 152, 0, 1, 
/* out0325_had-eta5-phi16*/	7, 61, 0, 5, 61, 1, 10, 102, 0, 3, 102, 2, 9, 103, 1, 1, 103, 2, 1, 151, 0, 4, 
/* out0326_had-eta6-phi16*/	7, 60, 0, 14, 60, 1, 4, 60, 2, 2, 61, 1, 1, 102, 2, 2, 150, 0, 3, 151, 0, 1, 
/* out0327_had-eta7-phi16*/	7, 49, 0, 1, 49, 1, 1, 59, 0, 5, 59, 2, 1, 60, 1, 9, 60, 2, 4, 150, 0, 3, 
/* out0328_had-eta8-phi16*/	5, 48, 0, 1, 49, 1, 1, 59, 0, 1, 59, 2, 13, 150, 0, 2, 
/* out0329_had-eta9-phi16*/	3, 48, 0, 6, 48, 1, 4, 59, 2, 2, 
/* out0330_had-eta10-phi16*/	3, 12, 0, 7, 48, 1, 8, 70, 2, 1, 
/* out0331_had-eta11-phi16*/	6, 12, 0, 6, 12, 1, 1, 12, 2, 14, 12, 3, 11, 12, 9, 1, 12, 10, 4, 
/* out0332_had-eta12-phi16*/	4, 12, 5, 4, 12, 6, 8, 12, 10, 12, 12, 11, 7, 
/* out0333_had-eta13-phi16*/	6, 11, 1, 3, 11, 7, 3, 12, 5, 7, 12, 11, 6, 16, 3, 3, 16, 9, 2, 
/* out0334_had-eta14-phi16*/	4, 11, 4, 3, 11, 7, 5, 16, 8, 3, 16, 9, 9, 
/* out0335_had-eta15-phi16*/	3, 5, 0, 5, 11, 4, 2, 16, 8, 10, 
/* out0336_had-eta16-phi16*/	3, 5, 0, 5, 5, 1, 8, 5, 2, 2, 
/* out0337_had-eta17-phi16*/	4, 5, 1, 1, 5, 2, 4, 5, 6, 6, 5, 7, 1, 
/* out0338_had-eta18-phi16*/	4, 5, 4, 1, 5, 5, 3, 5, 6, 6, 5, 7, 1, 
/* out0339_had-eta19-phi16*/	2, 5, 4, 2, 5, 5, 6, 
/* out0340_had-eta0-phi17*/	1, 153, 0, 2, 
/* out0341_had-eta1-phi17*/	1, 153, 0, 4, 
/* out0342_had-eta2-phi17*/	3, 104, 0, 1, 152, 0, 3, 153, 0, 2, 
/* out0343_had-eta3-phi17*/	5, 104, 0, 14, 104, 1, 15, 104, 2, 9, 116, 0, 1, 152, 0, 4, 
/* out0344_had-eta4-phi17*/	9, 102, 0, 1, 103, 0, 2, 103, 1, 8, 104, 1, 1, 104, 2, 1, 116, 0, 7, 116, 2, 14, 151, 0, 3, 152, 0, 1, 
/* out0345_had-eta5-phi17*/	5, 102, 0, 12, 102, 1, 11, 102, 2, 3, 116, 2, 2, 151, 0, 4, 
/* out0346_had-eta6-phi17*/	7, 60, 1, 2, 102, 1, 5, 102, 2, 2, 112, 0, 8, 112, 2, 5, 150, 0, 3, 151, 0, 1, 
/* out0347_had-eta7-phi17*/	4, 59, 0, 7, 60, 1, 1, 112, 2, 11, 150, 0, 3, 
/* out0348_had-eta8-phi17*/	3, 59, 0, 3, 59, 1, 13, 150, 0, 2, 
/* out0349_had-eta9-phi17*/	3, 59, 1, 3, 70, 0, 8, 70, 2, 3, 
/* out0350_had-eta10-phi17*/	2, 12, 0, 1, 70, 2, 11, 
/* out0351_had-eta11-phi17*/	6, 12, 0, 2, 12, 1, 15, 12, 2, 2, 12, 6, 2, 12, 7, 9, 70, 2, 1, 
/* out0352_had-eta12-phi17*/	4, 12, 4, 14, 12, 5, 3, 12, 6, 6, 12, 7, 7, 
/* out0353_had-eta13-phi17*/	5, 12, 4, 2, 12, 5, 2, 16, 0, 7, 16, 2, 1, 16, 3, 12, 
/* out0354_had-eta14-phi17*/	4, 16, 2, 6, 16, 3, 1, 16, 9, 5, 16, 10, 10, 
/* out0355_had-eta15-phi17*/	3, 16, 8, 3, 16, 10, 5, 16, 11, 10, 
/* out0356_had-eta16-phi17*/	3, 5, 1, 7, 5, 7, 1, 16, 11, 5, 
/* out0357_had-eta17-phi17*/	1, 5, 7, 11, 
/* out0358_had-eta18-phi17*/	2, 5, 4, 9, 5, 7, 2, 
/* out0359_had-eta19-phi17*/	1, 5, 4, 4, 
/* out0360_had-eta0-phi18*/	1, 157, 0, 2, 
/* out0361_had-eta1-phi18*/	1, 157, 0, 4, 
/* out0362_had-eta2-phi18*/	3, 117, 0, 1, 156, 0, 3, 157, 0, 2, 
/* out0363_had-eta3-phi18*/	5, 116, 0, 1, 117, 0, 14, 117, 1, 9, 117, 2, 15, 156, 0, 4, 
/* out0364_had-eta4-phi18*/	9, 113, 0, 1, 114, 0, 2, 114, 2, 8, 116, 0, 7, 116, 1, 14, 117, 1, 1, 117, 2, 1, 155, 0, 3, 156, 0, 1, 
/* out0365_had-eta5-phi18*/	5, 113, 0, 12, 113, 1, 3, 113, 2, 11, 116, 1, 2, 155, 0, 4, 
/* out0366_had-eta6-phi18*/	7, 72, 2, 2, 112, 0, 8, 112, 1, 5, 113, 1, 2, 113, 2, 5, 154, 0, 3, 155, 0, 1, 
/* out0367_had-eta7-phi18*/	4, 71, 0, 7, 72, 2, 1, 112, 1, 11, 154, 0, 3, 
/* out0368_had-eta8-phi18*/	3, 71, 0, 3, 71, 2, 13, 154, 0, 2, 
/* out0369_had-eta9-phi18*/	3, 70, 0, 8, 70, 1, 2, 71, 2, 3, 
/* out0370_had-eta10-phi18*/	2, 17, 0, 1, 70, 1, 10, 
/* out0371_had-eta11-phi18*/	6, 17, 0, 2, 17, 2, 2, 17, 3, 15, 17, 9, 9, 17, 10, 2, 70, 1, 2, 
/* out0372_had-eta12-phi18*/	4, 17, 8, 14, 17, 9, 7, 17, 10, 5, 17, 11, 3, 
/* out0373_had-eta13-phi18*/	5, 16, 0, 9, 16, 1, 11, 16, 2, 2, 17, 8, 2, 17, 11, 2, 
/* out0374_had-eta14-phi18*/	4, 16, 1, 1, 16, 2, 7, 16, 6, 10, 16, 7, 3, 
/* out0375_had-eta15-phi18*/	4, 16, 4, 1, 16, 5, 10, 16, 6, 6, 16, 10, 1, 
/* out0376_had-eta16-phi18*/	4, 16, 5, 6, 16, 11, 1, 21, 3, 7, 21, 9, 1, 
/* out0377_had-eta17-phi18*/	1, 21, 9, 11, 
/* out0378_had-eta18-phi18*/	2, 21, 8, 9, 21, 9, 2, 
/* out0379_had-eta19-phi18*/	1, 21, 8, 4, 
/* out0380_had-eta0-phi19*/	1, 157, 0, 2, 
/* out0381_had-eta1-phi19*/	1, 157, 0, 4, 
/* out0382_had-eta2-phi19*/	3, 115, 0, 3, 156, 0, 3, 157, 0, 2, 
/* out0383_had-eta3-phi19*/	7, 114, 0, 4, 115, 0, 10, 115, 1, 4, 115, 2, 16, 117, 0, 1, 117, 1, 6, 156, 0, 4, 
/* out0384_had-eta4-phi19*/	7, 73, 0, 1, 74, 2, 1, 114, 0, 10, 114, 1, 15, 114, 2, 7, 155, 0, 3, 156, 0, 1, 
/* out0385_had-eta5-phi19*/	7, 73, 0, 5, 73, 2, 10, 113, 0, 3, 113, 1, 9, 114, 1, 1, 114, 2, 1, 155, 0, 4, 
/* out0386_had-eta6-phi19*/	7, 72, 0, 14, 72, 1, 2, 72, 2, 4, 73, 2, 1, 113, 1, 2, 154, 0, 3, 155, 0, 1, 
/* out0387_had-eta7-phi19*/	7, 71, 0, 5, 71, 1, 1, 72, 1, 4, 72, 2, 9, 83, 0, 1, 83, 2, 1, 154, 0, 3, 
/* out0388_had-eta8-phi19*/	5, 71, 0, 1, 71, 1, 13, 82, 0, 1, 83, 2, 1, 154, 0, 2, 
/* out0389_had-eta9-phi19*/	4, 70, 1, 1, 71, 1, 2, 82, 0, 6, 82, 2, 4, 
/* out0390_had-eta10-phi19*/	3, 17, 0, 7, 70, 1, 1, 82, 2, 8, 
/* out0391_had-eta11-phi19*/	6, 17, 0, 6, 17, 1, 11, 17, 2, 14, 17, 3, 1, 17, 6, 4, 17, 7, 1, 
/* out0392_had-eta12-phi19*/	4, 17, 5, 7, 17, 6, 12, 17, 10, 9, 17, 11, 4, 
/* out0393_had-eta13-phi19*/	6, 16, 1, 4, 16, 7, 2, 17, 5, 6, 17, 11, 7, 22, 3, 3, 22, 9, 3, 
/* out0394_had-eta14-phi19*/	4, 16, 4, 4, 16, 7, 11, 22, 8, 3, 22, 9, 5, 
/* out0395_had-eta15-phi19*/	3, 16, 4, 11, 21, 0, 5, 22, 8, 2, 
/* out0396_had-eta16-phi19*/	3, 21, 0, 5, 21, 2, 2, 21, 3, 8, 
/* out0397_had-eta17-phi19*/	4, 21, 2, 4, 21, 3, 1, 21, 9, 1, 21, 10, 6, 
/* out0398_had-eta18-phi19*/	4, 21, 8, 1, 21, 9, 1, 21, 10, 6, 21, 11, 3, 
/* out0399_had-eta19-phi19*/	2, 21, 8, 2, 21, 11, 6, 
/* out0400_had-eta0-phi20*/	1, 161, 0, 2, 
/* out0401_had-eta1-phi20*/	1, 161, 0, 4, 
/* out0402_had-eta2-phi20*/	4, 75, 0, 5, 115, 0, 1, 160, 0, 3, 161, 0, 2, 
/* out0403_had-eta3-phi20*/	6, 74, 0, 10, 75, 0, 6, 75, 2, 15, 115, 0, 2, 115, 1, 12, 160, 0, 4, 
/* out0404_had-eta4-phi20*/	7, 73, 0, 4, 74, 0, 5, 74, 1, 9, 74, 2, 15, 85, 0, 1, 159, 0, 3, 160, 0, 1, 
/* out0405_had-eta5-phi20*/	6, 73, 0, 6, 73, 1, 15, 73, 2, 3, 84, 0, 1, 85, 2, 2, 159, 0, 4, 
/* out0406_had-eta6-phi20*/	8, 72, 0, 2, 72, 1, 6, 73, 1, 1, 73, 2, 2, 84, 0, 5, 84, 2, 8, 158, 0, 3, 159, 0, 1, 
/* out0407_had-eta7-phi20*/	5, 72, 1, 4, 83, 0, 12, 83, 2, 1, 84, 2, 2, 158, 0, 3, 
/* out0408_had-eta8-phi20*/	4, 82, 0, 1, 83, 1, 2, 83, 2, 13, 158, 0, 2, 
/* out0409_had-eta9-phi20*/	2, 82, 0, 8, 82, 1, 5, 
/* out0410_had-eta10-phi20*/	3, 23, 3, 2, 82, 1, 7, 82, 2, 4, 
/* out0411_had-eta11-phi20*/	6, 17, 1, 5, 17, 4, 1, 17, 7, 13, 23, 3, 5, 23, 8, 1, 23, 9, 11, 
/* out0412_had-eta12-phi20*/	5, 17, 4, 15, 17, 5, 2, 17, 7, 2, 22, 0, 5, 23, 8, 6, 
/* out0413_had-eta13-phi20*/	5, 17, 5, 1, 22, 0, 5, 22, 2, 5, 22, 3, 13, 22, 9, 1, 
/* out0414_had-eta14-phi20*/	5, 22, 2, 1, 22, 8, 3, 22, 9, 7, 22, 10, 10, 22, 11, 1, 
/* out0415_had-eta15-phi20*/	4, 21, 0, 4, 21, 1, 1, 22, 8, 8, 22, 11, 5, 
/* out0416_had-eta16-phi20*/	3, 21, 0, 2, 21, 1, 8, 21, 2, 5, 
/* out0417_had-eta17-phi20*/	3, 21, 2, 5, 21, 6, 7, 21, 10, 1, 
/* out0418_had-eta18-phi20*/	4, 21, 5, 2, 21, 6, 5, 21, 10, 3, 21, 11, 1, 
/* out0419_had-eta19-phi20*/	2, 21, 5, 4, 21, 11, 6, 
/* out0420_had-eta0-phi21*/	1, 161, 0, 2, 
/* out0421_had-eta1-phi21*/	1, 161, 0, 4, 
/* out0422_had-eta2-phi21*/	5, 75, 0, 4, 75, 1, 2, 87, 1, 5, 160, 0, 3, 161, 0, 2, 
/* out0423_had-eta3-phi21*/	10, 74, 0, 1, 74, 1, 1, 75, 0, 1, 75, 1, 14, 75, 2, 1, 86, 0, 14, 86, 1, 1, 86, 2, 4, 87, 1, 7, 160, 0, 4, 
/* out0424_had-eta4-phi21*/	7, 74, 1, 6, 85, 0, 13, 85, 1, 2, 86, 1, 1, 86, 2, 12, 159, 0, 3, 160, 0, 1, 
/* out0425_had-eta5-phi21*/	5, 84, 0, 4, 85, 0, 2, 85, 1, 8, 85, 2, 14, 159, 0, 4, 
/* out0426_had-eta6-phi21*/	6, 84, 0, 6, 84, 1, 13, 84, 2, 3, 95, 2, 1, 158, 0, 3, 159, 0, 1, 
/* out0427_had-eta7-phi21*/	7, 83, 0, 3, 83, 1, 4, 84, 1, 2, 84, 2, 3, 94, 0, 3, 94, 2, 4, 158, 0, 3, 
/* out0428_had-eta8-phi21*/	4, 83, 1, 10, 93, 0, 5, 94, 2, 1, 158, 0, 2, 
/* out0429_had-eta9-phi21*/	3, 82, 1, 2, 93, 0, 3, 93, 2, 8, 
/* out0430_had-eta10-phi21*/	6, 23, 0, 16, 23, 1, 4, 23, 2, 2, 23, 3, 5, 82, 1, 2, 93, 2, 2, 
/* out0431_had-eta11-phi21*/	5, 23, 2, 12, 23, 3, 4, 23, 6, 2, 23, 9, 5, 23, 10, 13, 
/* out0432_had-eta12-phi21*/	5, 22, 0, 4, 22, 1, 3, 23, 8, 9, 23, 10, 3, 23, 11, 12, 
/* out0433_had-eta13-phi21*/	5, 22, 0, 2, 22, 1, 11, 22, 2, 9, 22, 6, 3, 22, 7, 2, 
/* out0434_had-eta14-phi21*/	4, 22, 2, 1, 22, 5, 2, 22, 6, 12, 22, 10, 6, 
/* out0435_had-eta15-phi21*/	3, 21, 1, 1, 22, 5, 6, 22, 11, 10, 
/* out0436_had-eta16-phi21*/	2, 21, 1, 6, 21, 7, 8, 
/* out0437_had-eta17-phi21*/	3, 21, 4, 2, 21, 6, 3, 21, 7, 7, 
/* out0438_had-eta18-phi21*/	3, 21, 4, 5, 21, 5, 5, 21, 6, 1, 
/* out0439_had-eta19-phi21*/	1, 21, 5, 5, 
/* out0440_had-eta0-phi22*/	1, 165, 0, 2, 
/* out0441_had-eta1-phi22*/	1, 165, 0, 4, 
/* out0442_had-eta2-phi22*/	5, 87, 0, 5, 87, 1, 1, 97, 0, 1, 164, 0, 3, 165, 0, 2, 
/* out0443_had-eta3-phi22*/	7, 86, 0, 2, 86, 1, 7, 87, 0, 11, 87, 1, 3, 97, 0, 12, 97, 2, 12, 164, 0, 4, 
/* out0444_had-eta4-phi22*/	8, 85, 1, 2, 86, 1, 7, 96, 0, 14, 96, 1, 2, 96, 2, 8, 97, 2, 1, 163, 0, 3, 164, 0, 1, 
/* out0445_had-eta5-phi22*/	6, 85, 1, 4, 95, 0, 15, 95, 1, 2, 95, 2, 1, 96, 2, 7, 163, 0, 4, 
/* out0446_had-eta6-phi22*/	6, 84, 1, 1, 94, 0, 6, 95, 1, 3, 95, 2, 14, 162, 0, 3, 163, 0, 1, 
/* out0447_had-eta7-phi22*/	4, 94, 0, 7, 94, 1, 7, 94, 2, 5, 162, 0, 3, 
/* out0448_had-eta8-phi22*/	5, 93, 0, 6, 93, 1, 2, 94, 1, 2, 94, 2, 6, 162, 0, 2, 
/* out0449_had-eta9-phi22*/	3, 93, 0, 2, 93, 1, 9, 93, 2, 3, 
/* out0450_had-eta10-phi22*/	4, 23, 1, 12, 23, 7, 7, 93, 1, 2, 93, 2, 3, 
/* out0451_had-eta11-phi22*/	5, 23, 2, 2, 23, 4, 10, 23, 5, 3, 23, 6, 13, 23, 7, 9, 
/* out0452_had-eta12-phi22*/	5, 22, 1, 1, 23, 4, 2, 23, 5, 13, 23, 6, 1, 23, 11, 4, 
/* out0453_had-eta13-phi22*/	3, 22, 1, 1, 22, 4, 1, 22, 7, 12, 
/* out0454_had-eta14-phi22*/	4, 22, 4, 14, 22, 5, 3, 22, 6, 1, 22, 7, 2, 
/* out0455_had-eta15-phi22*/	2, 22, 4, 1, 22, 5, 5, 
/* out0456_had-eta16-phi22*/	0, 
/* out0457_had-eta17-phi22*/	2, 21, 4, 4, 21, 7, 1, 
/* out0458_had-eta18-phi22*/	1, 21, 4, 5, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	1, 165, 0, 2, 
/* out0461_had-eta1-phi23*/	1, 165, 0, 4, 
/* out0462_had-eta2-phi23*/	2, 164, 0, 3, 165, 0, 2, 
/* out0463_had-eta3-phi23*/	4, 97, 0, 3, 97, 1, 16, 97, 2, 2, 164, 0, 4, 
/* out0464_had-eta4-phi23*/	5, 96, 0, 2, 96, 1, 12, 97, 2, 1, 163, 0, 3, 164, 0, 1, 
/* out0465_had-eta5-phi23*/	5, 95, 0, 1, 95, 1, 5, 96, 1, 2, 96, 2, 1, 163, 0, 4, 
/* out0466_had-eta6-phi23*/	3, 95, 1, 6, 162, 0, 3, 163, 0, 1, 
/* out0467_had-eta7-phi23*/	2, 94, 1, 6, 162, 0, 3, 
/* out0468_had-eta8-phi23*/	2, 94, 1, 1, 162, 0, 2, 
/* out0469_had-eta9-phi23*/	1, 93, 1, 3, 
/* out0470_had-eta10-phi23*/	0, 
/* out0471_had-eta11-phi23*/	1, 23, 4, 4, 
/* out0472_had-eta12-phi23*/	0, 
/* out0473_had-eta13-phi23*/	0, 
/* out0474_had-eta14-phi23*/	0, 
/* out0475_had-eta15-phi23*/	0, 
/* out0476_had-eta16-phi23*/	0, 
/* out0477_had-eta17-phi23*/	0, 
/* out0478_had-eta18-phi23*/	0, 
/* out0479_had-eta19-phi23*/	0, 
};