parameter integer matrixH [0:8213] = {
/* num inputs = 198(in0-in197) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2577 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	2,142,0,16,142,1,3,
/* out0002_em-eta2-phi0*/	4,60,0,1,60,1,2,141,0,4,142,1,13,
/* out0003_em-eta3-phi0*/	6,59,1,1,60,0,15,60,1,1,60,2,2,141,0,12,141,1,6,
/* out0004_em-eta4-phi0*/	5,51,1,8,59,0,14,59,1,1,140,0,7,141,1,10,
/* out0005_em-eta5-phi0*/	10,50,1,2,51,0,16,51,1,8,51,2,16,58,0,8,58,1,1,59,0,1,59,2,1,140,0,9,140,1,8,
/* out0006_em-eta6-phi0*/	7,50,0,16,50,1,14,50,2,10,57,0,1,58,0,4,139,0,9,140,1,8,
/* out0007_em-eta7-phi0*/	5,49,1,7,50,2,6,57,0,6,139,0,7,139,1,10,
/* out0008_em-eta8-phi0*/	6,49,0,16,49,1,6,49,2,10,56,0,1,139,1,6,139,2,10,
/* out0009_em-eta9-phi0*/	5,48,1,8,49,2,3,56,0,3,138,0,8,139,2,6,
/* out0010_em-eta10-phi0*/	5,48,0,16,48,1,4,48,2,7,138,0,8,138,1,16,
/* out0011_em-eta11-phi0*/	8,6,3,5,7,2,16,7,3,13,10,5,2,11,5,2,48,2,5,104,0,4,104,1,9,
/* out0012_em-eta12-phi0*/	10,6,0,1,6,1,1,6,2,11,6,3,9,7,0,1,7,3,3,7,4,16,104,0,5,104,1,1,104,2,7,
/* out0013_em-eta13-phi0*/	8,6,1,10,6,2,5,7,0,15,7,1,7,103,0,3,103,1,7,104,0,7,104,2,2,
/* out0014_em-eta14-phi0*/	9,2,3,3,3,2,16,3,3,11,6,1,1,6,4,16,7,1,9,103,0,6,103,1,1,103,2,3,
/* out0015_em-eta15-phi0*/	8,2,2,7,2,3,4,3,3,5,3,4,5,102,0,1,102,1,2,103,0,7,103,2,4,
/* out0016_em-eta16-phi0*/	6,2,1,2,2,2,9,3,0,15,3,4,11,102,0,4,102,1,3,
/* out0017_em-eta17-phi0*/	5,2,1,1,3,0,1,3,1,11,102,0,4,102,2,1,
/* out0018_em-eta18-phi0*/	8,0,4,8,0,5,1,1,0,3,1,1,16,2,4,16,3,1,1,102,0,7,102,2,3,
/* out0019_em-eta19-phi0*/	6,0,0,16,0,2,15,0,3,9,1,0,9,1,3,4,1,5,4,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	2,142,2,3,142,3,16,
/* out0022_em-eta2-phi1*/	3,60,1,4,141,3,4,142,2,13,
/* out0023_em-eta3-phi1*/	7,59,1,2,60,1,9,60,2,14,70,0,10,70,1,2,141,2,6,141,3,12,
/* out0024_em-eta4-phi1*/	7,59,0,1,59,1,12,59,2,12,69,0,3,70,0,4,140,3,7,141,2,10,
/* out0025_em-eta5-phi1*/	7,58,0,3,58,1,15,58,2,4,59,2,3,69,0,3,140,2,8,140,3,9,
/* out0026_em-eta6-phi1*/	7,57,0,1,57,1,9,58,0,1,58,2,11,68,0,1,139,5,9,140,2,8,
/* out0027_em-eta7-phi1*/	5,57,0,7,57,1,4,57,2,7,139,4,10,139,5,7,
/* out0028_em-eta8-phi1*/	8,49,1,3,49,2,3,56,0,4,56,1,7,57,0,1,57,2,3,139,3,10,139,4,6,
/* out0029_em-eta9-phi1*/	6,48,1,3,56,0,8,56,1,1,56,2,4,138,3,8,139,3,6,
/* out0030_em-eta10-phi1*/	9,11,2,16,11,3,4,11,4,3,11,5,4,48,1,1,48,2,4,56,2,2,138,2,16,138,3,8,
/* out0031_em-eta11-phi1*/	6,10,5,13,11,0,7,11,4,6,11,5,10,100,2,10,104,1,6,
/* out0032_em-eta12-phi1*/	7,6,0,11,6,3,2,9,2,3,10,4,12,10,5,1,98,0,5,104,2,7,
/* out0033_em-eta13-phi1*/	6,6,0,4,6,1,4,9,2,7,9,5,10,98,0,4,103,1,6,
/* out0034_em-eta14-phi1*/	5,2,3,3,8,5,13,9,5,5,103,1,2,103,2,6,
/* out0035_em-eta15-phi1*/	6,2,0,8,2,3,6,8,4,3,97,0,1,102,1,2,103,2,3,
/* out0036_em-eta16-phi1*/	4,2,0,7,2,1,7,5,2,1,102,1,6,
/* out0037_em-eta17-phi1*/	5,2,1,6,3,1,1,5,5,5,102,1,1,102,2,5,
/* out0038_em-eta18-phi1*/	5,0,4,8,0,5,3,3,1,3,4,5,3,102,2,3,
/* out0039_em-eta19-phi1*/	6,0,2,1,0,3,5,0,5,8,1,0,4,1,3,10,1,5,10,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	2,147,0,16,147,1,3,
/* out0042_em-eta2-phi2*/	2,146,0,4,147,1,13,
/* out0043_em-eta3-phi2*/	8,70,0,2,70,1,14,70,2,8,79,0,2,80,1,1,80,2,11,146,0,12,146,1,6,
/* out0044_em-eta4-phi2*/	7,69,0,4,69,1,15,69,2,2,70,2,8,79,0,5,145,0,7,146,1,10,
/* out0045_em-eta5-phi2*/	7,58,2,1,68,0,1,68,1,7,69,0,6,69,2,12,145,0,9,145,1,8,
/* out0046_em-eta6-phi2*/	6,57,1,1,68,0,13,68,1,3,68,2,5,144,0,9,145,1,8,
/* out0047_em-eta7-phi2*/	8,57,1,2,57,2,5,67,0,7,67,1,3,68,0,1,68,2,1,144,0,7,144,1,10,
/* out0048_em-eta8-phi2*/	5,56,1,7,57,2,1,67,0,7,144,1,6,144,2,10,
/* out0049_em-eta9-phi2*/	5,56,1,1,56,2,9,66,0,3,143,0,8,144,2,6,
/* out0050_em-eta10-phi2*/	10,10,2,3,10,3,15,11,3,12,11,4,4,56,2,1,66,0,1,100,1,1,100,2,3,143,0,8,143,1,16,
/* out0051_em-eta11-phi2*/	10,10,0,1,10,1,6,10,2,13,10,3,1,11,0,9,11,1,2,11,4,3,98,1,3,100,1,13,100,2,3,
/* out0052_em-eta12-phi2*/	8,9,2,4,9,3,9,10,1,1,10,4,4,11,1,13,98,0,3,98,1,8,98,2,1,
/* out0053_em-eta13-phi2*/	7,8,2,2,9,2,2,9,3,5,9,4,14,9,5,1,98,0,4,98,2,6,
/* out0054_em-eta14-phi2*/	8,8,2,1,8,4,1,8,5,3,9,0,13,9,1,1,9,4,2,97,0,4,97,1,4,
/* out0055_em-eta15-phi2*/	5,2,0,1,5,2,3,8,4,12,9,1,2,97,0,7,
/* out0056_em-eta16-phi2*/	4,5,2,11,5,5,3,97,0,3,102,1,2,
/* out0057_em-eta17-phi2*/	6,4,5,1,5,0,1,5,4,3,5,5,8,96,1,2,102,2,3,
/* out0058_em-eta18-phi2*/	4,4,5,10,96,0,1,96,1,2,102,2,1,
/* out0059_em-eta19-phi2*/	5,0,3,2,0,5,4,1,3,2,1,5,2,4,4,4,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	2,147,2,3,147,3,16,
/* out0062_em-eta2-phi3*/	6,80,1,1,80,2,2,132,0,2,132,2,1,146,3,4,147,2,13,
/* out0063_em-eta3-phi3*/	9,79,0,1,79,1,15,79,2,1,80,1,14,80,2,3,132,0,1,132,2,12,146,2,6,146,3,12,
/* out0064_em-eta4-phi3*/	9,69,1,1,69,2,1,78,0,1,78,1,7,79,0,8,79,1,1,79,2,15,145,3,7,146,2,10,
/* out0065_em-eta5-phi3*/	7,68,1,3,69,2,1,78,0,15,78,1,3,78,2,5,145,2,8,145,3,9,
/* out0066_em-eta6-phi3*/	6,68,1,3,68,2,10,77,0,8,77,1,2,144,5,9,145,2,8,
/* out0067_em-eta7-phi3*/	6,67,0,1,67,1,13,67,2,3,77,0,2,144,4,10,144,5,7,
/* out0068_em-eta8-phi3*/	5,66,1,3,67,0,1,67,2,11,144,3,10,144,4,6,
/* out0069_em-eta9-phi3*/	5,66,0,6,66,1,6,66,2,1,143,3,8,144,3,6,
/* out0070_em-eta10-phi3*/	9,10,0,6,13,2,2,66,0,6,66,2,3,100,1,1,101,0,4,101,2,1,143,2,16,143,3,8,
/* out0071_em-eta11-phi3*/	8,10,0,9,10,1,6,13,2,11,13,5,9,100,1,1,101,0,4,101,1,1,101,2,12,
/* out0072_em-eta12-phi3*/	12,8,3,7,9,3,2,10,1,3,11,1,1,12,4,1,12,5,10,13,5,6,98,1,5,98,2,3,99,1,1,101,1,1,101,2,3,
/* out0073_em-eta13-phi3*/	7,8,0,6,8,1,1,8,2,8,8,3,9,97,1,1,98,2,6,99,1,4,
/* out0074_em-eta14-phi3*/	5,8,1,9,8,2,5,9,0,3,9,1,4,97,1,8,
/* out0075_em-eta15-phi3*/	6,5,2,1,5,3,7,9,1,9,97,0,1,97,1,1,97,2,6,
/* out0076_em-eta16-phi3*/	4,5,3,7,5,4,7,96,1,2,97,2,4,
/* out0077_em-eta17-phi3*/	4,4,2,1,5,0,5,5,4,6,96,1,5,
/* out0078_em-eta18-phi3*/	6,4,4,1,4,5,2,5,0,6,5,1,1,96,0,4,96,1,1,
/* out0079_em-eta19-phi3*/	1,4,4,9,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	2,152,0,16,152,1,3,
/* out0082_em-eta2-phi4*/	3,132,0,4,151,0,4,152,1,13,
/* out0083_em-eta3-phi4*/	9,131,0,1,131,1,9,132,0,9,132,1,16,132,2,3,133,1,1,133,2,6,151,0,12,151,1,6,
/* out0084_em-eta4-phi4*/	7,78,1,4,130,1,1,131,0,15,131,1,5,131,2,8,150,0,7,151,1,10,
/* out0085_em-eta5-phi4*/	7,77,1,2,78,1,2,78,2,11,130,0,10,130,1,2,150,0,9,150,1,8,
/* out0086_em-eta6-phi4*/	6,77,0,3,77,1,12,77,2,7,130,0,1,149,0,9,150,1,8,
/* out0087_em-eta7-phi4*/	7,67,2,1,76,0,2,76,1,6,77,0,3,77,2,6,149,0,7,149,1,10,
/* out0088_em-eta8-phi4*/	5,66,1,2,67,2,1,76,0,13,149,1,6,149,2,10,
/* out0089_em-eta9-phi4*/	5,66,1,5,66,2,6,76,0,1,148,0,8,149,2,6,
/* out0090_em-eta10-phi4*/	8,12,3,4,13,2,1,13,3,9,66,2,6,86,1,1,101,0,2,148,0,8,148,1,16,
/* out0091_em-eta11-phi4*/	9,12,2,8,12,3,2,13,0,1,13,2,2,13,3,7,13,4,15,13,5,1,101,0,6,101,1,11,
/* out0092_em-eta12-phi4*/	8,12,4,6,12,5,6,13,0,14,13,1,3,13,4,1,99,1,1,99,2,8,101,1,3,
/* out0093_em-eta13-phi4*/	7,8,0,8,12,4,8,14,5,4,15,5,3,99,0,1,99,1,7,99,2,1,
/* out0094_em-eta14-phi4*/	9,8,0,2,8,1,5,14,4,6,14,5,7,92,1,1,97,1,2,97,2,1,99,0,2,99,1,3,
/* out0095_em-eta15-phi4*/	6,4,3,6,5,3,2,8,1,1,14,4,7,92,1,3,97,2,4,
/* out0096_em-eta16-phi4*/	6,4,2,4,4,3,10,92,1,1,96,1,2,96,2,2,97,2,1,
/* out0097_em-eta17-phi4*/	5,4,1,1,4,2,10,5,0,1,96,1,2,96,2,3,
/* out0098_em-eta18-phi4*/	6,4,1,1,4,2,1,5,0,3,5,1,6,96,0,6,96,2,1,
/* out0099_em-eta19-phi4*/	3,4,4,2,5,1,4,96,0,2,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	2,152,2,3,152,3,16,
/* out0102_em-eta2-phi5*/	4,133,0,2,133,2,4,151,3,4,152,2,13,
/* out0103_em-eta3-phi5*/	7,120,1,4,131,1,1,133,0,14,133,1,15,133,2,6,151,2,6,151,3,12,
/* out0104_em-eta4-phi5*/	7,120,0,15,120,1,4,130,1,4,131,1,1,131,2,8,150,3,7,151,2,10,
/* out0105_em-eta5-phi5*/	5,130,0,4,130,1,9,130,2,14,150,2,8,150,3,9,
/* out0106_em-eta6-phi5*/	7,77,2,2,118,1,8,118,2,8,130,0,1,130,2,2,149,5,9,150,2,8,
/* out0107_em-eta7-phi5*/	6,76,1,9,76,2,1,77,2,1,118,1,8,149,4,10,149,5,7,
/* out0108_em-eta8-phi5*/	5,76,1,1,76,2,14,86,2,1,149,3,10,149,4,6,
/* out0109_em-eta9-phi5*/	5,76,2,1,86,1,5,86,2,7,148,3,8,149,3,6,
/* out0110_em-eta10-phi5*/	4,12,3,4,86,1,10,148,2,16,148,3,8,
/* out0111_em-eta11-phi5*/	7,12,0,16,12,1,5,12,2,6,12,3,6,94,0,9,94,1,1,94,2,10,
/* out0112_em-eta12-phi5*/	8,12,1,11,12,2,2,13,0,1,13,1,12,15,2,1,94,2,6,99,0,1,99,2,6,
/* out0113_em-eta13-phi5*/	8,12,4,1,13,1,1,14,5,1,15,2,6,15,4,4,15,5,13,99,0,9,99,2,1,
/* out0114_em-eta14-phi5*/	6,14,4,1,14,5,4,15,0,13,15,4,3,92,2,5,99,0,3,
/* out0115_em-eta15-phi5*/	5,14,4,2,15,0,3,15,1,12,92,1,5,92,2,2,
/* out0116_em-eta16-phi5*/	4,4,0,11,15,1,3,92,1,6,96,2,1,
/* out0117_em-eta17-phi5*/	3,4,0,5,4,1,7,96,2,5,
/* out0118_em-eta18-phi5*/	4,4,1,7,5,1,3,96,0,1,96,2,4,
/* out0119_em-eta19-phi5*/	2,5,1,2,96,0,2,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	2,157,0,16,157,1,3,
/* out0122_em-eta2-phi6*/	3,122,0,4,156,0,4,157,1,13,
/* out0123_em-eta3-phi6*/	7,120,1,4,121,2,1,122,0,12,122,1,10,122,2,16,156,0,12,156,1,6,
/* out0124_em-eta4-phi6*/	8,119,2,4,120,0,1,120,1,4,120,2,16,121,1,8,121,2,1,155,0,7,156,1,10,
/* out0125_em-eta5-phi6*/	5,119,0,4,119,1,14,119,2,9,155,0,9,155,1,8,
/* out0126_em-eta6-phi6*/	7,88,1,2,118,0,8,118,2,8,119,0,1,119,1,2,154,0,9,155,1,8,
/* out0127_em-eta7-phi6*/	6,87,1,1,87,2,9,88,1,1,118,0,8,154,0,7,154,1,10,
/* out0128_em-eta8-phi6*/	5,86,2,1,87,1,14,87,2,1,154,1,6,154,2,10,
/* out0129_em-eta9-phi6*/	5,86,0,4,86,2,7,87,1,1,153,0,8,154,2,6,
/* out0130_em-eta10-phi6*/	5,17,2,3,17,5,1,86,0,9,153,0,8,153,1,16,
/* out0131_em-eta11-phi6*/	7,16,5,13,17,0,4,17,4,2,17,5,14,86,0,1,94,0,7,94,1,10,
/* out0132_em-eta12-phi6*/	8,15,2,2,16,4,16,16,5,3,17,0,4,17,1,5,93,1,1,93,2,6,94,1,5,
/* out0133_em-eta13-phi6*/	6,15,2,7,15,3,12,15,4,5,17,1,1,93,1,9,93,2,1,
/* out0134_em-eta14-phi6*/	5,14,2,13,14,3,3,15,4,4,92,2,6,93,1,3,
/* out0135_em-eta15-phi6*/	6,14,0,1,14,1,13,14,2,3,15,1,1,92,0,5,92,2,2,
/* out0136_em-eta16-phi6*/	4,14,1,3,18,5,3,19,5,8,92,0,5,
/* out0137_em-eta17-phi6*/	3,18,4,1,18,5,11,105,1,4,
/* out0138_em-eta18-phi6*/	2,18,4,9,105,1,4,
/* out0139_em-eta19-phi6*/	2,18,4,2,105,0,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	2,157,2,3,157,3,16,
/* out0142_em-eta2-phi7*/	3,123,0,4,156,3,4,157,2,13,
/* out0143_em-eta3-phi7*/	8,121,0,1,121,2,9,122,1,6,123,0,10,123,1,5,123,2,16,156,2,6,156,3,12,
/* out0144_em-eta4-phi7*/	7,89,2,4,119,2,1,121,0,15,121,1,8,121,2,5,155,3,7,156,2,10,
/* out0145_em-eta5-phi7*/	7,88,2,2,89,1,11,89,2,2,119,0,10,119,2,2,155,2,8,155,3,9,
/* out0146_em-eta6-phi7*/	6,88,0,3,88,1,7,88,2,12,119,0,1,154,5,9,155,2,8,
/* out0147_em-eta7-phi7*/	7,87,0,2,87,2,6,88,0,3,88,1,6,99,1,1,154,4,10,154,5,7,
/* out0148_em-eta8-phi7*/	5,87,0,13,98,2,2,99,1,1,154,3,10,154,4,6,
/* out0149_em-eta9-phi7*/	6,86,0,1,87,0,1,98,1,6,98,2,5,153,3,8,154,3,6,
/* out0150_em-eta10-phi7*/	7,17,2,11,17,3,3,86,0,1,98,1,6,95,0,2,153,2,16,153,3,8,
/* out0151_em-eta11-phi7*/	10,16,2,8,16,3,1,17,0,2,17,2,2,17,3,8,17,4,14,17,5,1,95,0,8,95,1,1,95,2,11,
/* out0152_em-eta12-phi7*/	7,16,1,9,16,2,8,17,0,6,17,1,6,93,0,1,93,2,8,95,2,4,
/* out0153_em-eta13-phi7*/	9,14,3,5,15,3,4,16,1,4,17,1,4,20,5,4,21,5,3,93,0,7,93,1,1,93,2,1,
/* out0154_em-eta14-phi7*/	10,14,0,6,14,3,8,20,4,4,20,5,3,92,0,1,92,2,1,93,0,3,93,1,2,106,1,1,106,2,2,
/* out0155_em-eta15-phi7*/	5,14,0,9,19,2,8,20,4,1,92,0,3,106,1,4,
/* out0156_em-eta16-phi7*/	7,19,2,2,19,4,4,19,5,8,92,0,2,105,1,2,105,2,1,106,1,1,
/* out0157_em-eta17-phi7*/	5,18,5,2,19,0,8,19,4,2,105,1,4,105,2,1,
/* out0158_em-eta18-phi7*/	5,18,4,2,19,0,4,19,1,4,105,0,5,105,1,2,
/* out0159_em-eta19-phi7*/	3,18,4,2,19,1,5,105,0,2,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	2,162,0,16,162,1,3,
/* out0162_em-eta2-phi8*/	6,91,0,2,91,1,1,123,0,2,123,1,1,161,0,4,162,1,13,
/* out0163_em-eta3-phi8*/	8,90,0,1,90,1,1,90,2,15,91,0,3,91,1,14,123,1,10,161,0,12,161,1,6,
/* out0164_em-eta4-phi8*/	9,89,0,1,89,2,7,90,0,8,90,1,15,90,2,1,101,1,1,101,2,1,160,0,7,161,1,10,
/* out0165_em-eta5-phi8*/	7,89,0,15,89,1,5,89,2,3,100,2,3,101,1,1,160,0,9,160,1,8,
/* out0166_em-eta6-phi8*/	6,88,0,8,88,2,2,100,1,10,100,2,3,159,0,9,160,1,8,
/* out0167_em-eta7-phi8*/	6,88,0,2,99,0,1,99,1,3,99,2,13,159,0,7,159,1,10,
/* out0168_em-eta8-phi8*/	5,98,2,3,99,0,1,99,1,11,159,1,6,159,2,10,
/* out0169_em-eta9-phi8*/	5,98,0,6,98,1,1,98,2,6,158,0,8,159,2,6,
/* out0170_em-eta10-phi8*/	9,17,3,2,23,5,6,98,0,6,98,1,3,95,0,4,95,1,1,108,1,1,158,0,8,158,1,16,
/* out0171_em-eta11-phi8*/	9,16,0,3,16,3,15,17,3,3,22,4,3,22,5,11,23,5,1,95,0,2,95,1,12,108,1,1,
/* out0172_em-eta12-phi8*/	9,16,0,13,16,1,3,21,2,9,22,4,4,93,0,1,95,1,2,95,2,1,107,1,3,107,2,5,
/* out0173_em-eta13-phi8*/	8,20,5,3,21,0,2,21,2,2,21,4,6,21,5,13,93,0,4,106,2,1,107,1,6,
/* out0174_em-eta14-phi8*/	5,20,4,5,20,5,6,21,0,8,21,1,2,106,2,8,
/* out0175_em-eta15-phi8*/	7,19,2,5,19,3,3,20,4,6,21,1,3,106,0,1,106,1,6,106,2,1,
/* out0176_em-eta16-phi8*/	6,18,2,1,19,2,1,19,3,6,19,4,7,105,2,2,106,1,4,
/* out0177_em-eta17-phi8*/	4,18,2,8,19,0,2,19,4,3,105,2,6,
/* out0178_em-eta18-phi8*/	6,18,1,3,18,2,3,19,0,2,19,1,2,105,0,6,105,2,1,
/* out0179_em-eta19-phi8*/	2,18,1,3,19,1,5,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	2,162,2,3,162,3,16,
/* out0182_em-eta2-phi9*/	2,161,3,4,162,2,13,
/* out0183_em-eta3-phi9*/	8,90,0,2,91,0,11,91,1,1,102,0,2,102,1,8,102,2,14,161,2,6,161,3,12,
/* out0184_em-eta4-phi9*/	7,90,0,5,101,0,4,101,1,2,101,2,15,102,1,8,160,3,7,161,2,10,
/* out0185_em-eta5-phi9*/	7,100,0,1,100,2,7,101,0,6,101,1,12,110,1,1,160,2,8,160,3,9,
/* out0186_em-eta6-phi9*/	6,100,0,13,100,1,5,100,2,3,109,2,1,159,5,9,160,2,8,
/* out0187_em-eta7-phi9*/	8,99,0,7,99,2,3,100,0,1,100,1,1,109,1,5,109,2,2,159,4,10,159,5,7,
/* out0188_em-eta8-phi9*/	5,99,0,7,108,2,7,109,1,1,159,3,10,159,4,6,
/* out0189_em-eta9-phi9*/	5,98,0,3,108,1,9,108,2,1,158,3,8,159,3,6,
/* out0190_em-eta10-phi9*/	10,23,2,16,23,3,4,23,4,6,23,5,8,98,0,1,108,1,1,108,0,3,108,1,1,158,2,16,158,3,8,
/* out0191_em-eta11-phi9*/	10,22,2,2,22,4,2,22,5,5,23,0,16,23,1,2,23,4,8,23,5,1,107,2,3,108,0,3,108,1,13,
/* out0192_em-eta12-phi9*/	7,21,2,5,21,3,7,22,4,7,23,1,10,107,0,3,107,1,1,107,2,8,
/* out0193_em-eta13-phi9*/	6,20,2,6,20,3,2,21,3,7,21,4,10,107,0,4,107,1,6,
/* out0194_em-eta14-phi9*/	6,20,1,4,20,2,9,21,0,6,21,1,2,106,0,4,106,2,4,
/* out0195_em-eta15-phi9*/	4,19,3,3,20,1,5,21,1,9,106,0,7,
/* out0196_em-eta16-phi9*/	5,18,2,1,18,3,10,19,3,4,89,2,2,106,0,3,
/* out0197_em-eta17-phi9*/	5,18,0,4,18,2,3,18,3,5,89,1,3,105,2,3,
/* out0198_em-eta18-phi9*/	5,18,0,4,18,1,6,89,1,1,105,0,2,105,2,2,
/* out0199_em-eta19-phi9*/	5,18,1,4,24,3,3,24,5,1,25,3,2,25,5,2,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	2,167,0,16,167,1,3,
/* out0202_em-eta2-phi10*/	3,112,2,4,166,0,4,167,1,13,
/* out0203_em-eta3-phi10*/	7,102,0,10,102,2,2,111,2,2,112,1,14,112,2,9,166,0,12,166,1,6,
/* out0204_em-eta4-phi10*/	7,101,0,3,102,0,4,111,0,1,111,1,12,111,2,12,165,0,7,166,1,10,
/* out0205_em-eta5-phi10*/	7,101,0,3,110,0,3,110,1,4,110,2,15,111,1,3,165,0,9,165,1,8,
/* out0206_em-eta6-phi10*/	7,100,0,1,109,0,1,109,2,9,110,0,1,110,1,11,164,0,9,165,1,8,
/* out0207_em-eta7-phi10*/	5,109,0,7,109,1,7,109,2,4,164,0,7,164,1,10,
/* out0208_em-eta8-phi10*/	6,108,0,4,108,2,7,109,0,1,109,1,3,164,1,6,164,2,10,
/* out0209_em-eta9-phi10*/	5,108,0,8,108,1,4,108,2,1,163,0,8,164,2,6,
/* out0210_em-eta10-phi10*/	8,22,2,1,22,3,12,23,3,12,23,4,2,52,0,2,108,1,2,163,0,8,163,1,16,
/* out0211_em-eta11-phi10*/	6,22,0,12,22,1,7,22,2,13,22,3,4,91,2,6,108,0,10,
/* out0212_em-eta12-phi10*/	8,20,3,1,21,3,2,22,1,9,23,1,4,30,5,4,31,5,7,91,1,7,107,0,5,
/* out0213_em-eta13-phi10*/	6,20,0,4,20,3,13,30,4,2,30,5,5,90,2,6,107,0,4,
/* out0214_em-eta14-phi10*/	6,20,0,12,20,1,4,20,2,1,29,2,2,90,1,6,90,2,2,
/* out0215_em-eta15-phi10*/	7,20,1,3,28,5,1,29,2,1,29,5,12,89,2,2,90,1,3,106,0,1,
/* out0216_em-eta16-phi10*/	4,18,3,1,28,4,1,28,5,12,89,2,6,
/* out0217_em-eta17-phi10*/	4,18,0,5,28,4,6,89,1,5,89,2,1,
/* out0218_em-eta18-phi10*/	4,18,0,3,24,0,7,24,3,2,89,1,3,
/* out0219_em-eta19-phi10*/	5,24,2,1,24,3,9,24,5,5,25,3,9,25,5,9,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	2,167,2,3,167,3,16,
/* out0222_em-eta2-phi11*/	4,112,0,1,112,2,2,166,3,4,167,2,13,
/* out0223_em-eta3-phi11*/	6,111,2,1,112,0,15,112,1,2,112,2,1,166,2,6,166,3,12,
/* out0224_em-eta4-phi11*/	6,55,0,4,55,1,3,111,0,14,111,2,1,165,3,7,166,2,10,
/* out0225_em-eta5-phi11*/	9,54,1,1,55,0,12,55,2,4,110,0,8,110,2,1,111,0,1,111,1,1,165,2,8,165,3,9,
/* out0226_em-eta6-phi11*/	7,54,0,14,54,1,3,54,2,1,109,0,1,110,0,4,164,5,9,165,2,8,
/* out0227_em-eta7-phi11*/	7,53,0,3,53,1,3,54,0,2,54,2,3,109,0,6,164,4,10,164,5,7,
/* out0228_em-eta8-phi11*/	6,53,0,12,53,1,1,53,2,2,108,0,1,164,3,10,164,4,6,
/* out0229_em-eta9-phi11*/	7,52,0,4,52,1,3,53,0,1,53,2,2,108,0,3,163,3,8,164,3,6,
/* out0230_em-eta10-phi11*/	4,52,0,9,52,2,1,163,2,16,163,3,8,
/* out0231_em-eta11-phi11*/	7,22,0,4,31,2,13,31,3,2,52,0,1,52,2,3,91,0,4,91,2,9,
/* out0232_em-eta12-phi11*/	9,30,5,1,31,0,4,31,2,3,31,3,2,31,4,12,31,5,9,91,0,5,91,1,7,91,2,1,
/* out0233_em-eta13-phi11*/	7,30,4,8,30,5,6,31,0,8,31,1,3,90,0,2,90,2,7,91,1,2,
/* out0234_em-eta14-phi11*/	7,29,2,11,29,3,2,30,4,6,31,1,1,90,0,5,90,1,3,90,2,1,
/* out0235_em-eta15-phi11*/	7,29,2,2,29,3,1,29,4,11,29,5,4,89,2,2,90,0,1,90,1,4,
/* out0236_em-eta16-phi11*/	5,28,5,3,29,0,12,29,4,1,89,0,3,89,2,3,
/* out0237_em-eta17-phi11*/	4,28,4,8,29,1,3,89,0,4,89,1,1,
/* out0238_em-eta18-phi11*/	7,24,0,9,24,1,3,24,2,2,24,3,1,28,4,1,89,0,1,89,1,3,
/* out0239_em-eta19-phi11*/	6,24,2,8,24,3,1,24,5,8,25,0,4,25,3,5,25,5,5,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	2,172,0,16,172,1,3,
/* out0242_em-eta2-phi12*/	4,65,0,1,65,1,2,171,0,4,172,1,13,
/* out0243_em-eta3-phi12*/	6,64,1,1,65,0,15,65,1,1,65,2,2,171,0,12,171,1,6,
/* out0244_em-eta4-phi12*/	5,55,1,8,64,0,14,64,1,1,170,0,7,171,1,10,
/* out0245_em-eta5-phi12*/	9,54,1,1,55,1,5,55,2,12,63,0,8,63,1,1,64,0,1,64,2,1,170,0,9,170,1,8,
/* out0246_em-eta6-phi12*/	6,54,1,11,54,2,6,62,0,1,63,0,4,169,0,9,170,1,8,
/* out0247_em-eta7-phi12*/	5,53,1,7,54,2,6,62,0,6,169,0,7,169,1,10,
/* out0248_em-eta8-phi12*/	5,53,1,5,53,2,9,61,0,1,169,1,6,169,2,10,
/* out0249_em-eta9-phi12*/	5,52,1,8,53,2,3,61,0,3,168,0,8,169,2,6,
/* out0250_em-eta10-phi12*/	4,52,1,4,52,2,7,168,0,8,168,1,16,
/* out0251_em-eta11-phi12*/	8,30,3,5,31,3,10,36,5,2,37,5,2,52,2,4,88,0,11,88,2,1,91,0,3,
/* out0252_em-eta12-phi12*/	10,30,0,1,30,1,1,30,2,11,30,3,9,31,3,2,31,4,4,87,0,6,87,1,2,88,2,1,91,0,4,
/* out0253_em-eta13-phi12*/	6,30,1,10,30,2,5,31,0,4,31,1,6,87,0,8,90,0,2,
/* out0254_em-eta14-phi12*/	9,28,3,3,29,3,11,30,1,1,31,1,6,86,0,2,86,1,1,87,0,1,87,2,1,90,0,5,
/* out0255_em-eta15-phi12*/	6,28,2,7,28,3,4,29,3,2,29,4,4,86,0,6,90,0,1,
/* out0256_em-eta16-phi12*/	5,28,1,2,28,2,9,29,0,4,86,0,3,89,0,3,
/* out0257_em-eta17-phi12*/	4,28,1,1,29,1,11,85,0,2,89,0,4,
/* out0258_em-eta18-phi12*/	8,24,1,12,24,2,3,25,0,3,25,1,3,29,1,1,85,0,3,85,1,1,89,0,1,
/* out0259_em-eta19-phi12*/	5,24,2,2,24,4,5,24,5,2,25,0,9,25,1,2,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	2,172,2,3,172,3,16,
/* out0262_em-eta2-phi13*/	3,65,1,4,171,3,4,172,2,13,
/* out0263_em-eta3-phi13*/	7,64,1,2,65,1,9,65,2,14,75,0,10,75,1,2,171,2,6,171,3,12,
/* out0264_em-eta4-phi13*/	7,64,0,1,64,1,12,64,2,12,74,0,3,75,0,4,170,3,7,171,2,10,
/* out0265_em-eta5-phi13*/	7,63,0,3,63,1,15,63,2,4,64,2,3,74,0,3,170,2,8,170,3,9,
/* out0266_em-eta6-phi13*/	7,62,0,1,62,1,9,63,0,1,63,2,11,73,0,1,169,5,9,170,2,8,
/* out0267_em-eta7-phi13*/	5,62,0,7,62,1,4,62,2,7,169,4,10,169,5,7,
/* out0268_em-eta8-phi13*/	6,61,0,4,61,1,7,62,0,1,62,2,3,169,3,10,169,4,6,
/* out0269_em-eta9-phi13*/	5,61,0,8,61,1,1,61,2,4,168,3,8,169,3,6,
/* out0270_em-eta10-phi13*/	9,37,2,16,37,3,4,37,4,3,37,5,4,52,1,1,52,2,1,61,2,2,168,2,16,168,3,8,
/* out0271_em-eta11-phi13*/	7,36,5,13,37,0,7,37,4,6,37,5,10,84,0,1,88,0,5,88,2,13,
/* out0272_em-eta12-phi13*/	6,30,0,11,30,3,2,33,2,4,36,4,12,36,5,1,87,1,11,
/* out0273_em-eta13-phi13*/	6,30,0,4,30,1,4,33,2,6,33,5,10,87,0,1,87,2,8,
/* out0274_em-eta14-phi13*/	5,28,3,3,32,5,13,33,5,5,86,1,6,87,2,2,
/* out0275_em-eta15-phi13*/	6,28,0,8,28,3,6,32,4,3,86,0,3,86,1,2,86,2,1,
/* out0276_em-eta16-phi13*/	5,27,2,1,28,0,7,28,1,7,86,0,2,86,2,5,
/* out0277_em-eta17-phi13*/	4,27,5,5,28,1,6,29,1,1,85,0,6,
/* out0278_em-eta18-phi13*/	5,24,1,1,25,1,10,26,5,3,85,0,2,85,1,2,
/* out0279_em-eta19-phi13*/	2,24,4,8,25,1,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	2,177,0,16,177,1,3,
/* out0282_em-eta2-phi14*/	2,176,0,4,177,1,13,
/* out0283_em-eta3-phi14*/	8,75,0,2,75,1,14,75,2,8,84,0,2,85,0,11,85,2,1,176,0,12,176,1,6,
/* out0284_em-eta4-phi14*/	7,74,0,4,74,1,15,74,2,2,75,2,8,84,0,5,175,0,7,176,1,10,
/* out0285_em-eta5-phi14*/	7,63,2,1,73,0,1,73,1,7,74,0,6,74,2,12,175,0,9,175,1,8,
/* out0286_em-eta6-phi14*/	6,62,1,1,73,0,13,73,1,3,73,2,5,174,0,9,175,1,8,
/* out0287_em-eta7-phi14*/	8,62,1,2,62,2,5,72,0,7,72,1,3,73,0,1,73,2,1,174,0,7,174,1,10,
/* out0288_em-eta8-phi14*/	5,61,1,7,62,2,1,72,0,7,174,1,6,174,2,10,
/* out0289_em-eta9-phi14*/	5,61,1,1,61,2,9,71,0,3,173,0,8,174,2,6,
/* out0290_em-eta10-phi14*/	9,36,2,3,36,3,15,37,3,12,37,4,4,61,2,1,71,0,1,84,1,2,173,0,8,173,1,16,
/* out0291_em-eta11-phi14*/	10,36,0,1,36,1,6,36,2,13,36,3,1,37,0,9,37,1,2,37,4,3,84,0,9,84,1,5,88,2,1,
/* out0292_em-eta12-phi14*/	10,33,2,4,33,3,9,36,1,1,36,4,4,37,1,13,82,1,1,84,0,6,84,2,3,87,1,3,87,2,1,
/* out0293_em-eta13-phi14*/	7,32,2,2,33,2,2,33,3,5,33,4,14,33,5,1,82,0,6,87,2,4,
/* out0294_em-eta14-phi14*/	8,32,2,1,32,4,1,32,5,3,33,0,13,33,1,1,33,4,2,82,0,4,86,1,4,
/* out0295_em-eta15-phi14*/	6,27,2,3,28,0,1,32,4,12,33,1,2,86,1,3,86,2,4,
/* out0296_em-eta16-phi14*/	4,27,2,11,27,5,3,81,0,1,86,2,5,
/* out0297_em-eta17-phi14*/	6,26,5,1,27,0,1,27,4,3,27,5,8,85,0,3,85,1,4,
/* out0298_em-eta18-phi14*/	2,26,5,10,85,1,4,
/* out0299_em-eta19-phi14*/	2,24,4,3,26,4,4,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	2,177,2,3,177,3,16,
/* out0302_em-eta2-phi15*/	6,85,0,2,85,2,1,137,0,2,137,2,1,176,3,4,177,2,13,
/* out0303_em-eta3-phi15*/	9,84,0,1,84,1,15,84,2,1,85,0,3,85,2,14,137,0,1,137,2,12,176,2,6,176,3,12,
/* out0304_em-eta4-phi15*/	9,74,1,1,74,2,1,83,0,1,83,1,7,84,0,8,84,1,1,84,2,15,175,3,7,176,2,10,
/* out0305_em-eta5-phi15*/	7,73,1,3,74,2,1,83,0,15,83,1,3,83,2,5,175,2,8,175,3,9,
/* out0306_em-eta6-phi15*/	6,73,1,3,73,2,10,82,0,8,82,1,2,174,5,9,175,2,8,
/* out0307_em-eta7-phi15*/	6,72,0,1,72,1,13,72,2,3,82,0,2,174,4,10,174,5,7,
/* out0308_em-eta8-phi15*/	5,71,1,3,72,0,1,72,2,11,174,3,10,174,4,6,
/* out0309_em-eta9-phi15*/	5,71,0,6,71,1,6,71,2,1,173,3,8,174,3,6,
/* out0310_em-eta10-phi15*/	7,35,2,2,36,0,6,71,0,6,71,2,3,84,1,2,173,2,16,173,3,8,
/* out0311_em-eta11-phi15*/	6,35,2,11,35,5,9,36,0,9,36,1,6,84,1,7,84,2,6,
/* out0312_em-eta12-phi15*/	10,32,3,7,33,3,2,34,4,1,34,5,10,35,5,6,36,1,3,37,1,1,82,1,4,83,1,1,84,2,7,
/* out0313_em-eta13-phi15*/	7,32,0,6,32,1,1,32,2,8,32,3,9,82,0,3,82,1,7,82,2,1,
/* out0314_em-eta14-phi15*/	6,32,1,9,32,2,5,33,0,3,33,1,4,82,0,3,82,2,5,
/* out0315_em-eta15-phi15*/	7,27,2,1,27,3,7,33,1,9,81,0,3,81,1,3,82,2,1,86,2,1,
/* out0316_em-eta16-phi15*/	3,27,3,7,27,4,7,81,0,6,
/* out0317_em-eta17-phi15*/	5,26,2,1,27,0,5,27,4,6,81,0,3,85,1,3,
/* out0318_em-eta18-phi15*/	5,26,4,2,26,5,2,27,0,6,27,1,1,85,1,2,
/* out0319_em-eta19-phi15*/	1,26,4,8,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	2,182,0,16,182,1,3,
/* out0322_em-eta2-phi16*/	3,137,0,4,181,0,4,182,1,13,
/* out0323_em-eta3-phi16*/	9,135,0,1,135,1,9,136,1,1,136,2,6,137,0,9,137,1,16,137,2,3,181,0,12,181,1,6,
/* out0324_em-eta4-phi16*/	7,83,1,4,134,1,1,135,0,15,135,1,5,135,2,8,180,0,7,181,1,10,
/* out0325_em-eta5-phi16*/	7,82,1,2,83,1,2,83,2,11,134,0,10,134,1,2,180,0,9,180,1,8,
/* out0326_em-eta6-phi16*/	6,82,0,3,82,1,12,82,2,7,134,0,1,179,0,9,180,1,8,
/* out0327_em-eta7-phi16*/	7,72,2,1,81,0,2,81,1,6,82,0,3,82,2,6,179,0,7,179,1,10,
/* out0328_em-eta8-phi16*/	5,71,1,2,72,2,1,81,0,13,179,1,6,179,2,10,
/* out0329_em-eta9-phi16*/	5,71,1,5,71,2,6,81,0,1,178,0,8,179,2,6,
/* out0330_em-eta10-phi16*/	7,34,3,4,35,2,1,35,3,9,71,2,6,92,1,1,178,0,8,178,1,16,
/* out0331_em-eta11-phi16*/	9,34,2,8,34,3,2,35,0,1,35,2,2,35,3,7,35,4,15,35,5,1,83,1,4,83,2,8,
/* out0332_em-eta12-phi16*/	8,34,4,6,34,5,6,35,0,14,35,1,3,35,4,1,82,1,1,83,0,1,83,1,10,
/* out0333_em-eta13-phi16*/	9,32,0,8,34,4,8,38,5,4,39,5,3,79,0,1,82,1,3,82,2,4,83,0,1,83,1,1,
/* out0334_em-eta14-phi16*/	7,32,0,2,32,1,5,38,4,6,38,5,7,79,0,2,81,1,1,82,2,5,
/* out0335_em-eta15-phi16*/	5,26,3,6,27,3,2,32,1,1,38,4,7,81,1,7,
/* out0336_em-eta16-phi16*/	5,26,2,4,26,3,10,81,0,2,81,1,1,81,2,3,
/* out0337_em-eta17-phi16*/	5,26,1,1,26,2,10,27,0,1,81,0,1,81,2,3,
/* out0338_em-eta18-phi16*/	4,26,1,1,26,2,1,27,0,3,27,1,6,
/* out0339_em-eta19-phi16*/	2,26,4,2,27,1,4,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	2,182,2,3,182,3,16,
/* out0342_em-eta2-phi17*/	4,136,0,2,136,2,4,181,3,4,182,2,13,
/* out0343_em-eta3-phi17*/	7,128,1,4,135,1,1,136,0,14,136,1,15,136,2,6,181,2,6,181,3,12,
/* out0344_em-eta4-phi17*/	7,128,0,15,128,1,4,134,1,4,135,1,1,135,2,8,180,3,7,181,2,10,
/* out0345_em-eta5-phi17*/	5,134,0,4,134,1,9,134,2,14,180,2,8,180,3,9,
/* out0346_em-eta6-phi17*/	7,82,2,2,124,1,8,124,2,8,134,0,1,134,2,2,179,5,9,180,2,8,
/* out0347_em-eta7-phi17*/	6,81,1,9,81,2,1,82,2,1,124,1,8,179,4,10,179,5,7,
/* out0348_em-eta8-phi17*/	5,81,1,1,81,2,14,92,2,1,179,3,10,179,4,6,
/* out0349_em-eta9-phi17*/	5,81,2,1,92,1,5,92,2,7,178,3,8,179,3,6,
/* out0350_em-eta10-phi17*/	4,34,3,4,92,1,10,178,2,16,178,3,8,
/* out0351_em-eta11-phi17*/	6,34,0,16,34,1,5,34,2,6,34,3,6,83,0,2,83,2,8,
/* out0352_em-eta12-phi17*/	7,34,1,11,34,2,2,35,0,1,35,1,12,39,2,1,79,1,1,83,0,11,
/* out0353_em-eta13-phi17*/	9,34,4,1,35,1,1,38,5,1,39,2,6,39,4,4,39,5,13,79,0,3,79,1,7,83,0,1,
/* out0354_em-eta14-phi17*/	5,38,4,1,38,5,4,39,0,13,39,4,3,79,0,8,
/* out0355_em-eta15-phi17*/	6,38,4,2,39,0,2,39,1,12,79,0,2,81,1,4,81,2,1,
/* out0356_em-eta16-phi17*/	3,26,0,11,39,1,3,81,2,6,
/* out0357_em-eta17-phi17*/	3,26,0,5,26,1,7,81,2,3,
/* out0358_em-eta18-phi17*/	2,26,1,7,27,1,3,
/* out0359_em-eta19-phi17*/	1,27,1,2,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	2,187,0,16,187,1,3,
/* out0362_em-eta2-phi18*/	4,129,0,2,129,1,3,186,0,4,187,1,13,
/* out0363_em-eta3-phi18*/	7,126,2,1,128,1,4,129,0,14,129,1,8,129,2,15,186,0,12,186,1,6,
/* out0364_em-eta4-phi18*/	8,125,2,4,126,1,8,126,2,1,128,0,1,128,1,4,128,2,16,185,0,7,186,1,10,
/* out0365_em-eta5-phi18*/	5,125,0,4,125,1,14,125,2,9,185,0,9,185,1,8,
/* out0366_em-eta6-phi18*/	7,94,1,2,124,0,8,124,2,8,125,0,1,125,1,2,184,0,9,185,1,8,
/* out0367_em-eta7-phi18*/	6,93,1,1,93,2,9,94,1,1,124,0,8,184,0,7,184,1,10,
/* out0368_em-eta8-phi18*/	5,92,2,1,93,1,14,93,2,1,184,1,6,184,2,10,
/* out0369_em-eta9-phi18*/	5,92,0,4,92,2,7,93,1,1,183,0,8,184,2,6,
/* out0370_em-eta10-phi18*/	5,41,2,3,41,5,1,92,0,9,183,0,8,183,1,16,
/* out0371_em-eta11-phi18*/	7,40,5,13,41,0,4,41,4,2,41,5,14,92,0,1,80,0,2,80,1,8,
/* out0372_em-eta12-phi18*/	7,39,2,2,40,4,16,40,5,3,41,0,4,41,1,5,79,1,1,80,0,11,
/* out0373_em-eta13-phi18*/	7,39,2,7,39,3,12,39,4,5,41,1,1,79,1,7,79,2,2,80,0,1,
/* out0374_em-eta14-phi18*/	5,38,2,13,38,3,3,39,0,1,39,4,4,79,2,8,
/* out0375_em-eta15-phi18*/	7,38,0,1,38,1,13,38,2,3,39,1,1,76,1,1,76,2,4,79,2,2,
/* out0376_em-eta16-phi18*/	4,38,1,3,42,5,3,43,5,8,76,1,6,
/* out0377_em-eta17-phi18*/	3,42,4,1,42,5,11,76,1,3,
/* out0378_em-eta18-phi18*/	1,42,4,9,
/* out0379_em-eta19-phi18*/	1,42,4,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	2,187,2,3,187,3,16,
/* out0382_em-eta2-phi19*/	3,127,0,4,186,3,4,187,2,13,
/* out0383_em-eta3-phi19*/	9,126,0,1,126,2,9,127,0,10,127,1,5,127,2,16,129,1,5,129,2,1,186,2,6,186,3,12,
/* out0384_em-eta4-phi19*/	7,95,2,4,125,2,1,126,0,15,126,1,8,126,2,5,185,3,7,186,2,10,
/* out0385_em-eta5-phi19*/	7,94,2,2,95,1,11,95,2,2,125,0,10,125,2,2,185,2,8,185,3,9,
/* out0386_em-eta6-phi19*/	6,94,0,3,94,1,7,94,2,12,125,0,1,184,5,9,185,2,8,
/* out0387_em-eta7-phi19*/	7,93,0,2,93,2,6,94,0,3,94,1,6,104,1,1,184,4,10,184,5,7,
/* out0388_em-eta8-phi19*/	5,93,0,13,103,2,2,104,1,1,184,3,10,184,4,6,
/* out0389_em-eta9-phi19*/	6,92,0,1,93,0,1,103,1,6,103,2,5,183,3,8,184,3,6,
/* out0390_em-eta10-phi19*/	6,41,2,11,41,3,3,92,0,1,103,1,6,183,2,16,183,3,8,
/* out0391_em-eta11-phi19*/	9,40,2,8,40,3,1,41,0,2,41,2,2,41,3,8,41,4,14,41,5,1,80,1,8,80,2,4,
/* out0392_em-eta12-phi19*/	7,40,1,9,40,2,8,41,0,6,41,1,6,77,2,1,80,0,1,80,2,10,
/* out0393_em-eta13-phi19*/	11,38,3,5,39,3,4,40,1,4,41,1,4,44,5,4,45,5,3,77,1,4,77,2,3,79,2,2,80,0,1,80,2,1,
/* out0394_em-eta14-phi19*/	7,38,0,6,38,3,8,44,4,4,44,5,3,76,2,1,77,1,5,79,2,2,
/* out0395_em-eta15-phi19*/	4,38,0,9,43,2,8,44,4,1,76,2,7,
/* out0396_em-eta16-phi19*/	6,43,2,2,43,4,4,43,5,8,76,0,2,76,1,3,76,2,1,
/* out0397_em-eta17-phi19*/	5,42,5,2,43,0,8,43,4,2,76,0,1,76,1,3,
/* out0398_em-eta18-phi19*/	3,42,4,2,43,0,4,43,1,4,
/* out0399_em-eta19-phi19*/	2,42,4,2,43,1,5,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	2,192,0,16,192,1,3,
/* out0402_em-eta2-phi20*/	6,97,0,2,97,1,1,127,0,2,127,1,1,191,0,4,192,1,13,
/* out0403_em-eta3-phi20*/	8,96,0,1,96,1,1,96,2,15,97,0,3,97,1,14,127,1,10,191,0,12,191,1,6,
/* out0404_em-eta4-phi20*/	9,95,0,1,95,2,7,96,0,8,96,1,15,96,2,1,106,1,1,106,2,1,190,0,7,191,1,10,
/* out0405_em-eta5-phi20*/	7,95,0,15,95,1,5,95,2,3,105,2,3,106,1,1,190,0,9,190,1,8,
/* out0406_em-eta6-phi20*/	6,94,0,8,94,2,2,105,1,10,105,2,3,189,0,9,190,1,8,
/* out0407_em-eta7-phi20*/	6,94,0,2,104,0,1,104,1,3,104,2,13,189,0,7,189,1,10,
/* out0408_em-eta8-phi20*/	5,103,2,3,104,0,1,104,1,11,189,1,6,189,2,10,
/* out0409_em-eta9-phi20*/	5,103,0,6,103,1,1,103,2,6,188,0,8,189,2,6,
/* out0410_em-eta10-phi20*/	7,41,3,2,47,5,6,103,0,6,103,1,3,78,2,2,188,0,8,188,1,16,
/* out0411_em-eta11-phi20*/	8,40,0,3,40,3,15,41,3,3,46,4,3,46,5,11,47,5,1,78,1,6,78,2,7,
/* out0412_em-eta12-phi20*/	7,40,0,13,40,1,3,45,2,9,46,4,4,77,2,4,78,1,7,80,2,1,
/* out0413_em-eta13-phi20*/	8,44,5,3,45,0,2,45,2,2,45,4,6,45,5,13,77,0,3,77,1,1,77,2,7,
/* out0414_em-eta14-phi20*/	6,44,4,5,44,5,6,45,0,8,45,1,2,77,0,3,77,1,5,
/* out0415_em-eta15-phi20*/	8,43,2,5,43,3,3,44,4,6,45,1,3,73,1,1,76,0,3,76,2,3,77,1,1,
/* out0416_em-eta16-phi20*/	5,42,2,1,43,2,1,43,3,6,43,4,7,76,0,6,
/* out0417_em-eta17-phi20*/	5,42,2,8,43,0,2,43,4,3,72,1,3,76,0,3,
/* out0418_em-eta18-phi20*/	5,42,1,3,42,2,3,43,0,2,43,1,2,72,1,2,
/* out0419_em-eta19-phi20*/	2,42,1,3,43,1,5,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	2,192,2,3,192,3,16,
/* out0422_em-eta2-phi21*/	2,191,3,4,192,2,13,
/* out0423_em-eta3-phi21*/	8,96,0,2,97,0,11,97,1,1,107,0,2,107,1,8,107,2,14,191,2,6,191,3,12,
/* out0424_em-eta4-phi21*/	7,96,0,5,106,0,4,106,1,2,106,2,15,107,1,8,190,3,7,191,2,10,
/* out0425_em-eta5-phi21*/	7,105,0,1,105,2,7,106,0,6,106,1,12,115,1,1,190,2,8,190,3,9,
/* out0426_em-eta6-phi21*/	6,105,0,13,105,1,5,105,2,3,114,2,1,189,5,9,190,2,8,
/* out0427_em-eta7-phi21*/	8,104,0,7,104,2,3,105,0,1,105,1,1,114,1,5,114,2,2,189,4,10,189,5,7,
/* out0428_em-eta8-phi21*/	5,104,0,7,113,2,7,114,1,1,189,3,10,189,4,6,
/* out0429_em-eta9-phi21*/	5,103,0,3,113,1,9,113,2,1,188,3,8,189,3,6,
/* out0430_em-eta10-phi21*/	9,47,2,16,47,3,4,47,4,6,47,5,8,103,0,1,113,1,1,78,2,2,188,2,16,188,3,8,
/* out0431_em-eta11-phi21*/	10,46,2,2,46,4,2,46,5,5,47,0,16,47,1,2,47,4,8,47,5,1,75,1,1,78,0,9,78,2,5,
/* out0432_em-eta12-phi21*/	9,45,2,5,45,3,7,46,4,7,47,1,10,74,1,1,74,2,3,77,2,1,78,0,6,78,1,3,
/* out0433_em-eta13-phi21*/	6,44,2,6,44,3,2,45,3,7,45,4,10,74,1,4,77,0,6,
/* out0434_em-eta14-phi21*/	6,44,1,4,44,2,9,45,0,6,45,1,2,73,2,4,77,0,4,
/* out0435_em-eta15-phi21*/	5,43,3,3,44,1,5,45,1,9,73,1,4,73,2,3,
/* out0436_em-eta16-phi21*/	5,42,2,1,42,3,10,43,3,4,73,1,5,76,0,1,
/* out0437_em-eta17-phi21*/	5,42,0,4,42,2,3,42,3,5,72,1,4,72,2,3,
/* out0438_em-eta18-phi21*/	3,42,0,4,42,1,6,72,1,4,
/* out0439_em-eta19-phi21*/	1,42,1,4,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	2,197,0,16,197,1,3,
/* out0442_em-eta2-phi22*/	3,117,2,4,196,0,4,197,1,13,
/* out0443_em-eta3-phi22*/	7,107,0,10,107,2,2,116,2,2,117,1,14,117,2,9,196,0,12,196,1,6,
/* out0444_em-eta4-phi22*/	7,106,0,3,107,0,4,116,0,1,116,1,12,116,2,12,195,0,7,196,1,10,
/* out0445_em-eta5-phi22*/	7,106,0,3,115,0,3,115,1,4,115,2,15,116,1,3,195,0,9,195,1,8,
/* out0446_em-eta6-phi22*/	7,105,0,1,114,0,1,114,2,9,115,0,1,115,1,11,194,0,9,195,1,8,
/* out0447_em-eta7-phi22*/	5,114,0,7,114,1,7,114,2,4,194,0,7,194,1,10,
/* out0448_em-eta8-phi22*/	6,113,0,4,113,2,7,114,0,1,114,1,3,194,1,6,194,2,10,
/* out0449_em-eta9-phi22*/	5,113,0,8,113,1,4,113,2,1,193,0,8,194,2,6,
/* out0450_em-eta10-phi22*/	7,46,2,1,46,3,12,47,3,12,47,4,2,113,1,2,193,0,8,193,1,16,
/* out0451_em-eta11-phi22*/	7,46,0,12,46,1,7,46,2,13,46,3,4,75,0,5,75,1,13,78,0,1,
/* out0452_em-eta12-phi22*/	5,44,3,1,45,3,2,46,1,9,47,1,4,74,2,11,
/* out0453_em-eta13-phi22*/	4,44,0,4,44,3,13,74,0,1,74,1,8,
/* out0454_em-eta14-phi22*/	5,44,0,12,44,1,4,44,2,1,73,2,6,74,1,2,
/* out0455_em-eta15-phi22*/	4,44,1,3,73,0,3,73,1,1,73,2,2,
/* out0456_em-eta16-phi22*/	3,42,3,1,73,0,2,73,1,5,
/* out0457_em-eta17-phi22*/	2,42,0,5,72,2,6,
/* out0458_em-eta18-phi22*/	3,42,0,3,72,1,2,72,2,2,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	2,197,2,3,197,3,16,
/* out0462_em-eta2-phi23*/	4,117,0,1,117,2,2,196,3,4,197,2,13,
/* out0463_em-eta3-phi23*/	6,116,2,1,117,0,15,117,1,2,117,2,1,196,2,6,196,3,12,
/* out0464_em-eta4-phi23*/	4,116,0,14,116,2,1,195,3,7,196,2,10,
/* out0465_em-eta5-phi23*/	6,115,0,8,115,2,1,116,0,1,116,1,1,195,2,8,195,3,9,
/* out0466_em-eta6-phi23*/	4,114,0,1,115,0,4,194,5,9,195,2,8,
/* out0467_em-eta7-phi23*/	3,114,0,6,194,4,10,194,5,7,
/* out0468_em-eta8-phi23*/	3,113,0,1,194,3,10,194,4,6,
/* out0469_em-eta9-phi23*/	3,113,0,3,193,3,8,194,3,6,
/* out0470_em-eta10-phi23*/	2,193,2,16,193,3,8,
/* out0471_em-eta11-phi23*/	3,46,0,4,75,0,11,75,1,1,
/* out0472_em-eta12-phi23*/	3,74,0,6,74,2,2,75,1,1,
/* out0473_em-eta13-phi23*/	1,74,0,8,
/* out0474_em-eta14-phi23*/	4,73,0,2,73,2,1,74,0,1,74,1,1,
/* out0475_em-eta15-phi23*/	1,73,0,6,
/* out0476_em-eta16-phi23*/	1,73,0,3,
/* out0477_em-eta17-phi23*/	1,72,2,2,
/* out0478_em-eta18-phi23*/	2,72,1,1,72,2,3,
/* out0479_em-eta19-phi23*/	0
};