parameter integer matrixH [0:5531] = {
/* num inputs = 140(in0-in139) */
/* num outputs = 600(out0-out599) */
//* max inputs per outputs = 8 */
//* total number of input in adders 1643 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	0,
/* out0006_em-eta6-phi0*/	0,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	0,
/* out0010_em-eta10-phi0*/	0,
/* out0011_em-eta11-phi0*/	0,
/* out0012_em-eta12-phi0*/	0,
/* out0013_em-eta13-phi0*/	0,
/* out0014_em-eta14-phi0*/	0,
/* out0015_em-eta15-phi0*/	0,
/* out0016_em-eta16-phi0*/	0,
/* out0017_em-eta17-phi0*/	0,
/* out0018_em-eta18-phi0*/	0,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	0,
/* out0026_em-eta6-phi1*/	0,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	0,
/* out0029_em-eta9-phi1*/	0,
/* out0030_em-eta10-phi1*/	0,
/* out0031_em-eta11-phi1*/	0,
/* out0032_em-eta12-phi1*/	0,
/* out0033_em-eta13-phi1*/	0,
/* out0034_em-eta14-phi1*/	0,
/* out0035_em-eta15-phi1*/	0,
/* out0036_em-eta16-phi1*/	0,
/* out0037_em-eta17-phi1*/	0,
/* out0038_em-eta18-phi1*/	0,
/* out0039_em-eta19-phi1*/	0,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	0,
/* out0046_em-eta6-phi2*/	0,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	0,
/* out0049_em-eta9-phi2*/	0,
/* out0050_em-eta10-phi2*/	0,
/* out0051_em-eta11-phi2*/	0,
/* out0052_em-eta12-phi2*/	0,
/* out0053_em-eta13-phi2*/	0,
/* out0054_em-eta14-phi2*/	0,
/* out0055_em-eta15-phi2*/	0,
/* out0056_em-eta16-phi2*/	0,
/* out0057_em-eta17-phi2*/	0,
/* out0058_em-eta18-phi2*/	0,
/* out0059_em-eta19-phi2*/	0,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	0,
/* out0065_em-eta5-phi3*/	0,
/* out0066_em-eta6-phi3*/	0,
/* out0067_em-eta7-phi3*/	0,
/* out0068_em-eta8-phi3*/	0,
/* out0069_em-eta9-phi3*/	0,
/* out0070_em-eta10-phi3*/	0,
/* out0071_em-eta11-phi3*/	0,
/* out0072_em-eta12-phi3*/	0,
/* out0073_em-eta13-phi3*/	0,
/* out0074_em-eta14-phi3*/	0,
/* out0075_em-eta15-phi3*/	0,
/* out0076_em-eta16-phi3*/	0,
/* out0077_em-eta17-phi3*/	0,
/* out0078_em-eta18-phi3*/	0,
/* out0079_em-eta19-phi3*/	0,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	4,60,0,1,60,1,3,77,0,10,77,1,15,
/* out0084_em-eta4-phi4*/	2,59,1,7,60,0,7,
/* out0085_em-eta5-phi4*/	3,59,0,15,59,1,6,59,2,5,
/* out0086_em-eta6-phi4*/	3,40,0,3,59,0,1,59,2,1,
/* out0087_em-eta7-phi4*/	2,39,0,2,39,1,10,
/* out0088_em-eta8-phi4*/	1,39,0,13,
/* out0089_em-eta9-phi4*/	1,39,0,1,
/* out0090_em-eta10-phi4*/	2,19,0,1,19,1,5,
/* out0091_em-eta11-phi4*/	4,19,0,15,19,1,5,19,2,7,19,3,7,
/* out0092_em-eta12-phi4*/	4,19,2,2,19,3,9,20,3,13,20,4,2,
/* out0093_em-eta13-phi4*/	1,20,2,1,
/* out0094_em-eta14-phi4*/	0,
/* out0095_em-eta15-phi4*/	0,
/* out0096_em-eta16-phi4*/	2,0,1,4,1,1,8,
/* out0097_em-eta17-phi4*/	2,0,0,1,0,1,11,
/* out0098_em-eta18-phi4*/	1,0,0,10,
/* out0099_em-eta19-phi4*/	1,0,0,2,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	3,61,1,1,61,2,10,77,0,1,
/* out0103_em-eta3-phi5*/	8,42,0,1,60,1,11,60,2,2,61,0,5,61,1,15,61,2,4,77,0,5,77,1,1,
/* out0104_em-eta4-phi5*/	5,41,0,6,59,1,2,60,0,8,60,1,2,60,2,14,
/* out0105_em-eta5-phi5*/	6,40,0,2,40,1,2,41,0,8,41,2,3,59,1,1,59,2,10,
/* out0106_em-eta6-phi5*/	3,40,0,11,40,1,6,40,2,6,
/* out0107_em-eta7-phi5*/	4,22,0,2,39,1,6,39,2,4,40,2,7,
/* out0108_em-eta8-phi5*/	3,21,1,2,22,0,1,39,2,12,
/* out0109_em-eta9-phi5*/	2,21,0,7,21,1,5,
/* out0110_em-eta10-phi5*/	4,19,1,4,19,4,2,20,1,11,21,0,5,
/* out0111_em-eta11-phi5*/	7,19,1,2,19,2,7,19,4,2,19,5,1,20,0,16,20,1,5,20,4,2,
/* out0112_em-eta12-phi5*/	4,20,2,8,20,3,3,20,4,12,20,5,6,
/* out0113_em-eta13-phi5*/	2,2,0,9,20,2,7,
/* out0114_em-eta14-phi5*/	2,2,0,1,2,3,5,
/* out0115_em-eta15-phi5*/	2,0,4,8,2,3,1,
/* out0116_em-eta16-phi5*/	3,0,4,2,1,0,4,1,1,8,
/* out0117_em-eta17-phi5*/	3,0,1,1,0,2,8,1,0,3,
/* out0118_em-eta18-phi5*/	3,0,0,2,0,2,4,0,3,4,
/* out0119_em-eta19-phi5*/	2,0,0,1,0,3,5,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	3,43,1,7,61,0,3,61,2,2,
/* out0123_em-eta3-phi6*/	5,42,0,10,42,1,11,43,0,7,43,1,6,61,0,8,
/* out0124_em-eta4-phi6*/	6,24,0,1,24,1,1,41,0,1,41,1,10,42,0,5,42,2,14,
/* out0125_em-eta5-phi6*/	6,23,1,5,24,0,1,40,1,1,41,0,1,41,1,6,41,2,13,
/* out0126_em-eta6-phi6*/	5,22,1,1,23,0,10,23,1,1,40,1,7,40,2,2,
/* out0127_em-eta7-phi6*/	4,22,0,11,22,1,5,22,2,1,40,2,1,
/* out0128_em-eta8-phi6*/	3,21,1,4,22,0,2,22,2,8,
/* out0129_em-eta9-phi6*/	3,21,0,1,21,1,5,21,2,7,
/* out0130_em-eta10-phi6*/	5,4,1,1,5,1,7,19,4,3,21,0,3,21,2,5,
/* out0131_em-eta11-phi6*/	4,4,0,4,4,1,10,19,4,9,19,5,11,
/* out0132_em-eta12-phi6*/	5,2,1,8,3,1,2,4,0,3,19,5,4,20,5,10,
/* out0133_em-eta13-phi6*/	4,2,0,6,2,1,8,2,2,9,2,3,1,
/* out0134_em-eta14-phi6*/	4,2,2,5,2,3,9,3,3,5,3,4,3,
/* out0135_em-eta15-phi6*/	3,0,4,5,0,5,3,3,3,8,
/* out0136_em-eta16-phi6*/	4,0,4,1,0,5,6,1,0,6,1,4,1,
/* out0137_em-eta17-phi6*/	3,0,2,2,1,0,3,1,4,8,
/* out0138_em-eta18-phi6*/	4,0,2,2,0,3,2,1,3,3,1,4,3,
/* out0139_em-eta19-phi6*/	2,0,3,5,1,3,3,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	1,43,1,1,
/* out0143_em-eta3-phi7*/	6,25,0,11,25,1,14,25,2,2,42,1,4,43,0,9,43,1,2,
/* out0144_em-eta4-phi7*/	6,24,0,4,24,1,15,24,2,5,25,0,5,42,1,1,42,2,2,
/* out0145_em-eta5-phi7*/	5,8,0,1,23,1,8,23,2,2,24,0,10,24,2,4,
/* out0146_em-eta6-phi7*/	4,7,1,2,23,0,6,23,1,2,23,2,13,
/* out0147_em-eta7-phi7*/	4,7,0,5,7,1,1,22,1,10,22,2,1,
/* out0148_em-eta8-phi7*/	3,6,0,8,6,1,1,22,2,6,
/* out0149_em-eta9-phi7*/	3,6,0,7,6,2,3,21,2,3,
/* out0150_em-eta10-phi7*/	5,4,4,16,4,5,4,5,0,9,5,1,8,21,2,1,
/* out0151_em-eta11-phi7*/	7,4,0,3,4,1,5,4,2,16,4,3,3,5,0,5,5,1,1,5,4,2,
/* out0152_em-eta12-phi7*/	4,2,4,4,3,1,10,4,0,6,4,3,9,
/* out0153_em-eta13-phi7*/	5,2,2,2,2,4,2,2,5,1,3,0,15,3,1,4,
/* out0154_em-eta14-phi7*/	5,3,0,1,3,2,1,3,3,2,3,4,13,3,5,3,
/* out0155_em-eta15-phi7*/	4,0,5,3,3,2,12,3,3,1,26,1,1,
/* out0156_em-eta16-phi7*/	3,0,5,4,1,4,1,1,5,10,
/* out0157_em-eta17-phi7*/	3,1,2,4,1,4,3,1,5,5,
/* out0158_em-eta18-phi7*/	2,1,2,4,1,3,6,
/* out0159_em-eta19-phi7*/	5,1,3,4,11,1,1,11,5,2,12,1,2,12,5,4,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	1,10,2,5,
/* out0163_em-eta3-phi8*/	5,9,1,5,10,1,14,10,2,10,25,1,2,25,2,12,
/* out0164_em-eta4-phi8*/	5,9,0,15,9,1,9,9,2,1,24,2,5,25,2,2,
/* out0165_em-eta5-phi8*/	4,8,0,6,8,1,15,8,2,3,24,2,2,
/* out0166_em-eta6-phi8*/	5,7,1,10,7,2,1,8,0,9,8,2,1,23,2,1,
/* out0167_em-eta7-phi8*/	3,7,0,9,7,1,3,7,2,7,
/* out0168_em-eta8-phi8*/	3,6,0,1,6,1,12,7,0,2,
/* out0169_em-eta9-phi8*/	2,6,1,1,6,2,10,
/* out0170_em-eta10-phi8*/	7,4,5,12,5,0,2,5,2,1,5,4,2,5,5,13,6,2,1,62,0,2,
/* out0171_em-eta11-phi8*/	4,5,2,11,5,3,8,5,4,12,5,5,3,
/* out0172_em-eta12-phi8*/	5,2,4,4,4,3,4,5,3,8,44,0,12,44,1,1,
/* out0173_em-eta13-phi8*/	4,2,4,6,2,5,11,44,0,3,44,3,4,
/* out0174_em-eta14-phi8*/	3,2,5,4,3,5,13,26,4,3,
/* out0175_em-eta15-phi8*/	4,3,2,3,26,1,1,26,4,1,27,1,13,
/* out0176_em-eta16-phi8*/	3,1,5,1,26,0,1,26,1,12,
/* out0177_em-eta17-phi8*/	2,1,2,5,26,0,6,
/* out0178_em-eta18-phi8*/	3,1,2,3,12,2,8,12,5,2,
/* out0179_em-eta19-phi8*/	5,11,1,5,11,5,10,12,1,10,12,4,1,12,5,9,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	5,9,1,1,9,2,1,10,1,2,10,2,1,114,1,1,
/* out0184_em-eta4-phi9*/	6,9,0,1,9,1,1,9,2,14,102,1,10,114,1,2,114,2,3,
/* out0185_em-eta5-phi9*/	6,8,1,1,8,2,9,90,0,1,90,1,2,102,0,12,102,1,2,
/* out0186_em-eta6-phi9*/	5,7,2,2,8,2,3,90,0,14,90,1,2,90,2,1,
/* out0187_em-eta7-phi9*/	5,7,2,6,78,0,5,78,1,4,90,0,1,90,2,3,
/* out0188_em-eta8-phi9*/	3,6,1,1,78,0,11,78,2,3,
/* out0189_em-eta9-phi9*/	5,6,1,1,6,2,2,62,0,5,62,1,4,78,2,1,
/* out0190_em-eta10-phi9*/	2,62,0,8,62,2,2,
/* out0191_em-eta11-phi9*/	5,5,2,4,44,1,6,45,1,11,62,0,1,62,2,2,
/* out0192_em-eta12-phi9*/	6,44,0,1,44,1,9,44,2,12,44,3,1,45,0,4,45,1,1,
/* out0193_em-eta13-phi9*/	4,44,2,4,44,3,10,45,3,7,45,4,4,
/* out0194_em-eta14-phi9*/	4,26,4,11,26,5,3,44,3,1,45,3,5,
/* out0195_em-eta15-phi9*/	4,26,4,1,26,5,1,27,0,12,27,1,3,
/* out0196_em-eta16-phi9*/	2,26,1,2,26,2,12,
/* out0197_em-eta17-phi9*/	2,26,0,8,26,3,4,
/* out0198_em-eta18-phi9*/	5,12,2,8,12,3,4,12,4,2,12,5,1,26,0,1,
/* out0199_em-eta19-phi9*/	5,11,1,8,11,2,4,11,5,4,12,1,4,12,4,9,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	5,114,1,13,114,2,3,115,1,2,125,1,2,125,2,12,
/* out0204_em-eta4-phi10*/	5,102,1,4,102,2,6,114,2,10,115,0,8,115,1,7,
/* out0205_em-eta5-phi10*/	5,90,1,3,102,0,4,102,2,10,103,0,3,103,1,7,
/* out0206_em-eta6-phi10*/	4,90,1,9,90,2,8,91,1,2,103,0,3,
/* out0207_em-eta7-phi10*/	4,78,1,8,90,2,4,91,0,3,91,1,3,
/* out0208_em-eta8-phi10*/	3,78,1,4,78,2,10,79,0,1,
/* out0209_em-eta9-phi10*/	3,62,1,8,78,2,2,79,0,2,
/* out0210_em-eta10-phi10*/	2,62,1,3,62,2,8,
/* out0211_em-eta11-phi10*/	4,44,4,14,45,1,3,62,2,3,63,0,4,
/* out0212_em-eta12-phi10*/	6,44,4,2,44,5,8,45,0,12,45,1,1,45,4,5,45,5,2,
/* out0213_em-eta13-phi10*/	4,45,2,8,45,3,3,45,4,7,45,5,5,
/* out0214_em-eta14-phi10*/	4,26,5,11,27,5,4,45,2,5,45,3,1,
/* out0215_em-eta15-phi10*/	4,26,5,1,27,0,4,27,4,8,27,5,4,
/* out0216_em-eta16-phi10*/	3,26,2,4,27,3,2,27,4,8,
/* out0217_em-eta17-phi10*/	2,26,3,10,27,3,2,
/* out0218_em-eta18-phi10*/	5,11,2,2,11,3,3,12,3,11,12,4,3,26,3,1,
/* out0219_em-eta19-phi10*/	5,11,0,5,11,1,2,11,2,10,11,3,2,12,4,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	6,115,1,3,115,2,1,125,1,14,125,2,4,126,0,12,126,1,2,
/* out0224_em-eta4-phi11*/	5,115,0,8,115,1,4,115,2,15,116,0,5,126,0,2,
/* out0225_em-eta5-phi11*/	4,103,0,3,103,1,9,103,2,12,116,0,2,
/* out0226_em-eta6-phi11*/	4,91,1,8,91,2,3,103,0,7,103,2,2,
/* out0227_em-eta7-phi11*/	3,91,0,10,91,1,3,91,2,5,
/* out0228_em-eta8-phi11*/	3,79,0,5,79,1,8,91,0,3,
/* out0229_em-eta9-phi11*/	2,79,0,8,79,2,5,
/* out0230_em-eta10-phi11*/	8,62,1,1,62,2,1,63,0,1,63,1,13,63,2,2,64,0,2,64,1,12,79,2,1,
/* out0231_em-eta11-phi11*/	4,63,0,11,63,1,3,63,2,12,63,3,8,
/* out0232_em-eta12-phi11*/	6,44,5,8,45,5,4,46,1,2,47,1,2,63,3,8,64,3,4,
/* out0233_em-eta13-phi11*/	4,45,2,3,45,5,5,46,0,5,46,1,12,
/* out0234_em-eta14-phi11*/	4,27,5,3,46,0,11,46,2,1,46,3,5,
/* out0235_em-eta15-phi11*/	3,27,2,9,27,5,5,46,3,3,
/* out0236_em-eta16-phi11*/	3,27,2,6,27,3,6,28,1,1,
/* out0237_em-eta17-phi11*/	3,26,3,1,27,3,6,28,0,5,
/* out0238_em-eta18-phi11*/	3,11,3,10,12,3,1,28,0,3,
/* out0239_em-eta19-phi11*/	2,11,0,8,11,3,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	1,134,2,1,
/* out0243_em-eta3-phi12*/	6,126,0,2,126,1,14,126,2,11,127,0,4,134,0,9,134,2,2,
/* out0244_em-eta4-phi12*/	5,116,0,5,116,1,15,116,2,4,126,2,5,127,0,3,
/* out0245_em-eta5-phi12*/	5,103,2,2,104,1,10,104,2,1,116,0,4,116,2,10,
/* out0246_em-eta6-phi12*/	4,91,2,2,104,0,13,104,1,6,104,2,1,
/* out0247_em-eta7-phi12*/	3,91,2,6,92,0,1,92,1,10,
/* out0248_em-eta8-phi12*/	3,79,1,8,79,2,1,92,0,6,
/* out0249_em-eta9-phi12*/	2,79,2,9,80,1,3,
/* out0250_em-eta10-phi12*/	5,63,4,16,63,5,8,64,0,9,64,1,4,80,0,1,
/* out0251_em-eta11-phi12*/	7,63,2,2,63,5,1,64,0,5,64,2,3,64,3,3,64,4,16,64,5,5,
/* out0252_em-eta12-phi12*/	4,46,4,5,47,1,8,64,2,6,64,3,9,
/* out0253_em-eta13-phi12*/	4,46,1,2,46,2,7,47,0,10,47,1,6,
/* out0254_em-eta14-phi12*/	4,46,2,8,46,3,4,47,3,2,47,4,6,
/* out0255_em-eta15-phi12*/	4,27,2,1,29,1,3,46,3,4,47,3,8,
/* out0256_em-eta16-phi12*/	3,28,1,10,28,2,1,29,1,4,
/* out0257_em-eta17-phi12*/	3,28,0,4,28,1,5,28,2,3,
/* out0258_em-eta18-phi12*/	2,28,0,4,28,3,6,
/* out0259_em-eta19-phi12*/	2,11,0,3,28,3,4,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	3,134,2,7,135,0,3,135,1,3,
/* out0263_em-eta3-phi13*/	6,127,0,3,127,1,16,127,2,3,134,0,7,134,2,6,135,0,10,
/* out0264_em-eta4-phi13*/	6,116,1,1,116,2,1,117,0,2,117,1,9,127,0,6,127,2,12,
/* out0265_em-eta5-phi13*/	6,104,2,5,105,1,1,116,2,1,117,0,14,117,1,1,117,2,5,
/* out0266_em-eta6-phi13*/	5,92,1,1,104,0,3,104,2,9,105,0,9,105,1,1,
/* out0267_em-eta7-phi13*/	4,92,0,1,92,1,5,92,2,11,105,0,1,
/* out0268_em-eta8-phi13*/	3,80,1,4,92,0,8,92,2,2,
/* out0269_em-eta9-phi13*/	3,80,0,3,80,1,9,80,2,1,
/* out0270_em-eta10-phi13*/	4,63,5,7,64,5,1,66,1,3,80,0,8,
/* out0271_em-eta11-phi13*/	5,64,2,4,64,5,10,65,0,4,65,1,15,66,1,2,
/* out0272_em-eta12-phi13*/	5,46,4,10,46,5,1,64,2,3,65,0,12,65,3,3,
/* out0273_em-eta13-phi13*/	5,46,4,1,46,5,12,47,0,6,47,4,3,47,5,3,
/* out0274_em-eta14-phi13*/	4,47,2,5,47,3,3,47,4,7,47,5,5,
/* out0275_em-eta15-phi13*/	4,28,4,5,29,1,3,47,2,6,47,3,3,
/* out0276_em-eta16-phi13*/	4,28,2,1,28,4,1,29,0,6,29,1,6,
/* out0277_em-eta17-phi13*/	3,28,2,8,29,0,3,29,4,2,
/* out0278_em-eta18-phi13*/	4,28,2,3,28,3,3,29,3,2,29,4,2,
/* out0279_em-eta19-phi13*/	2,28,3,3,29,3,5,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	2,135,1,10,135,2,1,
/* out0283_em-eta3-phi14*/	7,127,2,1,128,1,9,128,2,4,135,0,3,135,1,3,135,2,15,136,0,7,
/* out0284_em-eta4-phi14*/	5,117,1,5,118,1,2,128,0,14,128,1,7,128,2,3,
/* out0285_em-eta5-phi14*/	5,105,1,4,117,1,1,117,2,11,118,0,10,118,1,1,
/* out0286_em-eta6-phi14*/	3,105,0,4,105,1,10,105,2,8,
/* out0287_em-eta7-phi14*/	4,92,2,2,93,1,10,105,0,2,105,2,5,
/* out0288_em-eta8-phi14*/	4,80,2,2,92,2,1,93,0,7,93,1,4,
/* out0289_em-eta9-phi14*/	3,80,2,11,81,1,1,93,0,1,
/* out0290_em-eta10-phi14*/	5,65,4,12,66,1,5,80,0,4,80,2,2,81,1,1,
/* out0291_em-eta11-phi14*/	7,65,1,1,65,2,9,65,4,1,65,5,1,66,0,13,66,1,6,66,4,3,
/* out0292_em-eta12-phi14*/	4,65,2,7,65,3,10,66,3,6,66,4,5,
/* out0293_em-eta13-phi14*/	6,46,5,3,47,5,5,48,1,5,49,1,4,65,3,3,66,3,4,
/* out0294_em-eta14-phi14*/	4,47,2,4,47,5,3,48,0,7,48,1,7,
/* out0295_em-eta15-phi14*/	3,28,4,8,47,2,1,48,0,8,
/* out0296_em-eta16-phi14*/	3,28,4,2,28,5,8,29,0,4,
/* out0297_em-eta17-phi14*/	3,29,0,3,29,4,8,29,5,1,
/* out0298_em-eta18-phi14*/	3,29,2,2,29,3,4,29,4,4,
/* out0299_em-eta19-phi14*/	2,29,2,1,29,3,5,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	4,128,2,3,129,1,7,136,0,9,136,2,16,
/* out0304_em-eta4-phi15*/	5,118,1,7,128,0,2,128,2,6,129,0,8,129,1,9,
/* out0305_em-eta5-phi15*/	4,106,1,1,118,0,5,118,1,6,118,2,15,
/* out0306_em-eta6-phi15*/	5,105,2,3,106,0,10,106,1,7,118,0,1,118,2,1,
/* out0307_em-eta7-phi15*/	3,93,1,2,93,2,10,106,0,6,
/* out0308_em-eta8-phi15*/	3,81,1,1,93,0,8,93,2,6,
/* out0309_em-eta9-phi15*/	1,81,1,12,
/* out0310_em-eta10-phi15*/	4,65,4,3,65,5,3,81,0,8,81,1,1,
/* out0311_em-eta11-phi15*/	4,65,5,12,66,0,3,66,4,5,66,5,14,
/* out0312_em-eta12-phi15*/	5,48,4,3,66,2,16,66,3,5,66,4,3,66,5,2,
/* out0313_em-eta13-phi15*/	5,48,1,1,48,4,5,49,0,5,49,1,12,66,3,1,
/* out0314_em-eta14-phi15*/	3,48,1,3,48,2,14,49,0,3,
/* out0315_em-eta15-phi15*/	3,48,0,1,48,2,2,48,3,13,
/* out0316_em-eta16-phi15*/	3,28,5,8,29,5,4,48,3,3,
/* out0317_em-eta17-phi15*/	2,29,2,1,29,5,11,
/* out0318_em-eta18-phi15*/	1,29,2,10,
/* out0319_em-eta19-phi15*/	1,29,2,2,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	4,129,2,7,130,1,3,137,1,9,137,2,16,
/* out0324_em-eta4-phi16*/	6,119,1,4,119,2,3,129,0,8,129,2,9,130,0,2,130,1,6,
/* out0325_em-eta5-phi16*/	4,106,1,1,119,0,11,119,1,12,119,2,3,
/* out0326_em-eta6-phi16*/	4,106,1,7,106,2,10,107,0,3,119,0,1,
/* out0327_em-eta7-phi16*/	3,94,0,2,94,1,10,106,2,6,
/* out0328_em-eta8-phi16*/	2,81,2,1,94,0,13,
/* out0329_em-eta9-phi16*/	2,81,2,12,94,0,1,
/* out0330_em-eta10-phi16*/	4,67,4,1,67,5,5,81,0,8,81,2,1,
/* out0331_em-eta11-phi16*/	4,67,4,15,67,5,5,68,0,7,68,1,7,
/* out0332_em-eta12-phi16*/	5,48,4,3,67,1,13,67,2,2,68,0,2,68,1,9,
/* out0333_em-eta13-phi16*/	5,48,4,5,48,5,12,49,0,5,49,5,1,67,0,1,
/* out0334_em-eta14-phi16*/	3,49,0,3,49,4,14,49,5,3,
/* out0335_em-eta15-phi16*/	3,49,2,1,49,3,13,49,4,2,
/* out0336_em-eta16-phi16*/	2,30,4,11,49,3,3,
/* out0337_em-eta17-phi16*/	2,30,4,5,31,1,7,
/* out0338_em-eta18-phi16*/	2,30,1,3,31,1,7,
/* out0339_em-eta19-phi16*/	1,30,1,2,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	2,138,0,2,138,1,5,
/* out0343_em-eta3-phi17*/	7,130,1,4,130,2,9,131,0,1,137,1,7,138,0,14,138,1,3,138,2,12,
/* out0344_em-eta4-phi17*/	5,119,2,2,120,1,6,130,0,14,130,1,3,130,2,7,
/* out0345_em-eta5-phi17*/	5,107,1,4,119,0,4,119,2,8,120,0,3,120,1,8,
/* out0346_em-eta6-phi17*/	3,107,0,8,107,1,10,107,2,4,
/* out0347_em-eta7-phi17*/	5,94,1,6,94,2,4,95,0,1,107,0,5,107,2,2,
/* out0348_em-eta8-phi17*/	3,82,1,2,94,2,12,95,0,1,
/* out0349_em-eta9-phi17*/	2,81,2,1,82,1,11,
/* out0350_em-eta10-phi17*/	6,67,5,4,68,2,2,68,5,11,81,2,1,82,0,4,82,1,2,
/* out0351_em-eta11-phi17*/	7,67,2,2,67,5,2,68,0,7,68,2,2,68,3,1,68,4,16,68,5,5,
/* out0352_em-eta12-phi17*/	4,67,0,8,67,1,3,67,2,12,67,3,6,
/* out0353_em-eta13-phi17*/	4,48,5,4,49,5,5,50,4,9,67,0,7,
/* out0354_em-eta14-phi17*/	4,49,2,7,49,5,7,50,4,1,51,1,5,
/* out0355_em-eta15-phi17*/	4,30,5,7,31,5,2,49,2,8,51,1,1,
/* out0356_em-eta16-phi17*/	2,30,5,9,31,0,4,
/* out0357_em-eta17-phi17*/	3,30,2,1,31,0,10,31,1,1,
/* out0358_em-eta18-phi17*/	4,30,1,6,30,2,3,31,0,1,31,1,1,
/* out0359_em-eta19-phi17*/	2,30,0,3,30,1,4,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	2,138,1,4,139,0,7,
/* out0363_em-eta3-phi18*/	7,131,0,3,131,1,16,131,2,3,138,1,4,138,2,4,139,0,6,139,2,7,
/* out0364_em-eta4-phi18*/	5,120,1,1,120,2,10,121,1,3,131,0,12,131,2,6,
/* out0365_em-eta5-phi18*/	6,107,1,1,108,1,5,120,0,13,120,1,1,120,2,6,121,1,1,
/* out0366_em-eta6-phi18*/	5,95,1,1,107,1,1,107,2,9,108,0,3,108,1,9,
/* out0367_em-eta7-phi18*/	4,95,0,4,95,1,12,95,2,1,107,2,1,
/* out0368_em-eta8-phi18*/	3,82,2,4,95,0,10,95,2,1,
/* out0369_em-eta9-phi18*/	3,82,0,3,82,1,1,82,2,9,
/* out0370_em-eta10-phi18*/	3,68,2,3,69,4,7,82,0,8,
/* out0371_em-eta11-phi18*/	4,68,2,9,68,3,11,69,4,7,70,1,7,
/* out0372_em-eta12-phi18*/	6,50,5,8,51,5,2,67,3,10,68,3,4,69,1,1,70,1,2,
/* out0373_em-eta13-phi18*/	4,50,4,6,50,5,8,51,0,9,51,1,1,
/* out0374_em-eta14-phi18*/	4,50,1,5,50,2,3,51,0,5,51,1,9,
/* out0375_em-eta15-phi18*/	3,31,2,1,31,5,7,50,1,8,
/* out0376_em-eta16-phi18*/	2,31,4,7,31,5,7,
/* out0377_em-eta17-phi18*/	3,30,2,5,31,0,1,31,4,6,
/* out0378_em-eta18-phi18*/	4,30,0,1,30,1,1,30,2,6,30,3,2,
/* out0379_em-eta19-phi18*/	1,30,0,8,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	1,139,0,1,
/* out0383_em-eta3-phi19*/	6,131,2,4,132,0,11,132,1,14,132,2,2,139,0,2,139,2,9,
/* out0384_em-eta4-phi19*/	5,121,0,2,121,1,10,121,2,12,131,2,3,132,0,5,
/* out0385_em-eta5-phi19*/	5,108,1,1,108,2,10,109,1,2,121,0,12,121,1,2,
/* out0386_em-eta6-phi19*/	4,96,1,2,108,0,13,108,1,1,108,2,6,
/* out0387_em-eta7-phi19*/	3,95,1,3,95,2,8,96,1,6,
/* out0388_em-eta8-phi19*/	3,83,1,8,83,2,1,95,2,6,
/* out0389_em-eta9-phi19*/	3,82,2,3,83,0,3,83,1,7,
/* out0390_em-eta10-phi19*/	6,69,4,1,69,5,16,70,0,4,70,4,5,70,5,12,82,0,1,
/* out0391_em-eta11-phi19*/	6,69,1,4,69,2,9,69,4,1,70,0,12,70,1,7,70,4,2,
/* out0392_em-eta12-phi19*/	4,51,2,4,51,5,10,69,0,4,69,1,11,
/* out0393_em-eta13-phi19*/	5,51,0,2,51,2,2,51,3,1,51,4,15,51,5,4,
/* out0394_em-eta14-phi19*/	5,50,0,1,50,1,2,50,2,13,50,3,3,51,4,1,
/* out0395_em-eta15-phi19*/	4,31,2,4,32,1,1,50,0,12,50,1,1,
/* out0396_em-eta16-phi19*/	3,31,2,10,31,3,3,31,4,1,
/* out0397_em-eta17-phi19*/	4,30,2,1,30,3,1,31,3,8,31,4,2,
/* out0398_em-eta18-phi19*/	1,30,3,10,
/* out0399_em-eta19-phi19*/	2,13,4,3,30,0,4,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	2,133,0,3,133,2,1,
/* out0403_em-eta3-phi20*/	6,122,1,1,122,2,3,132,1,2,132,2,12,133,0,13,133,2,12,
/* out0404_em-eta4-phi20*/	5,121,2,4,122,0,8,122,1,15,122,2,4,132,2,2,
/* out0405_em-eta5-phi20*/	4,109,0,3,109,1,12,109,2,9,121,0,2,
/* out0406_em-eta6-phi20*/	4,96,1,3,96,2,8,109,0,7,109,1,2,
/* out0407_em-eta7-phi20*/	3,96,0,10,96,1,5,96,2,3,
/* out0408_em-eta8-phi20*/	3,83,1,1,83,2,12,96,0,3,
/* out0409_em-eta9-phi20*/	2,83,0,10,83,2,1,
/* out0410_em-eta10-phi20*/	6,70,2,16,70,3,6,70,4,4,70,5,4,71,1,2,83,0,1,
/* out0411_em-eta11-phi20*/	4,69,2,7,69,3,14,70,3,8,70,4,5,
/* out0412_em-eta12-phi20*/	4,51,2,4,52,1,4,53,1,8,69,0,12,
/* out0413_em-eta13-phi20*/	4,51,2,6,51,3,11,52,0,3,52,1,5,
/* out0414_em-eta14-phi20*/	3,32,4,3,50,3,13,51,3,4,
/* out0415_em-eta15-phi20*/	4,32,1,1,32,4,1,33,1,13,50,0,3,
/* out0416_em-eta16-phi20*/	3,31,2,1,32,0,1,32,1,12,
/* out0417_em-eta17-phi20*/	2,31,3,5,32,0,6,
/* out0418_em-eta18-phi20*/	3,13,5,10,14,5,1,30,3,3,
/* out0419_em-eta19-phi20*/	2,13,4,8,13,5,1,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	2,122,2,2,133,2,3,
/* out0424_em-eta4-phi21*/	4,110,1,10,122,0,8,122,2,7,123,2,5,
/* out0425_em-eta5-phi21*/	5,97,1,3,109,0,3,109,2,7,110,0,12,110,1,2,
/* out0426_em-eta6-phi21*/	4,96,2,2,97,0,8,97,1,9,109,0,3,
/* out0427_em-eta7-phi21*/	5,84,1,5,84,2,4,96,0,3,96,2,3,97,0,4,
/* out0428_em-eta8-phi21*/	3,83,2,1,84,0,3,84,1,11,
/* out0429_em-eta9-phi21*/	5,71,1,5,71,2,4,83,0,2,83,2,1,84,0,1,
/* out0430_em-eta10-phi21*/	2,71,0,2,71,1,8,
/* out0431_em-eta11-phi21*/	6,52,4,14,52,5,3,69,3,2,70,3,2,71,0,2,71,1,1,
/* out0432_em-eta12-phi21*/	6,52,1,2,52,2,5,52,4,2,52,5,1,53,0,12,53,1,8,
/* out0433_em-eta13-phi21*/	4,52,0,8,52,1,5,52,2,7,52,3,3,
/* out0434_em-eta14-phi21*/	4,32,4,11,32,5,3,52,0,5,52,3,1,
/* out0435_em-eta15-phi21*/	4,32,4,1,32,5,1,33,0,12,33,1,3,
/* out0436_em-eta16-phi21*/	2,32,1,2,32,2,12,
/* out0437_em-eta17-phi21*/	2,32,0,8,32,3,4,
/* out0438_em-eta18-phi21*/	5,13,5,3,14,0,2,14,4,3,14,5,11,32,0,1,
/* out0439_em-eta19-phi21*/	5,13,4,5,13,5,2,14,0,10,14,1,2,14,4,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	2,124,0,2,124,1,4,
/* out0443_em-eta3-phi22*/	7,111,1,1,111,2,1,123,1,12,123,2,5,124,0,14,124,1,2,124,2,3,
/* out0444_em-eta4-phi22*/	7,110,1,4,110,2,6,111,0,1,111,1,14,111,2,1,123,1,4,123,2,6,
/* out0445_em-eta5-phi22*/	6,97,1,2,97,2,1,98,1,9,98,2,1,110,0,4,110,2,10,
/* out0446_em-eta6-phi22*/	5,85,1,2,97,0,1,97,1,2,97,2,14,98,1,3,
/* out0447_em-eta7-phi22*/	4,84,2,8,85,1,6,97,0,3,97,2,1,
/* out0448_em-eta8-phi22*/	3,72,1,1,84,0,10,84,2,4,
/* out0449_em-eta9-phi22*/	3,71,2,8,72,1,2,84,0,2,
/* out0450_em-eta10-phi22*/	2,71,0,8,71,2,3,
/* out0451_em-eta11-phi22*/	4,52,5,11,53,5,6,54,4,4,71,0,3,
/* out0452_em-eta12-phi22*/	6,52,5,1,53,0,4,53,2,1,53,3,1,53,4,12,53,5,9,
/* out0453_em-eta13-phi22*/	4,52,2,4,52,3,7,53,3,10,53,4,4,
/* out0454_em-eta14-phi22*/	4,32,5,11,33,5,4,52,3,5,53,3,1,
/* out0455_em-eta15-phi22*/	4,32,5,1,33,0,4,33,4,8,33,5,4,
/* out0456_em-eta16-phi22*/	3,32,2,4,33,3,2,33,4,8,
/* out0457_em-eta17-phi22*/	2,32,3,10,33,3,2,
/* out0458_em-eta18-phi22*/	5,14,2,8,14,3,1,14,4,2,14,5,4,32,3,1,
/* out0459_em-eta19-phi22*/	5,13,1,4,13,3,4,14,0,4,14,1,8,14,4,9,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	1,124,1,2,
/* out0463_em-eta3-phi23*/	5,111,2,5,112,1,12,112,2,2,124,1,8,124,2,13,
/* out0464_em-eta4-phi23*/	5,99,1,4,111,0,15,111,1,1,111,2,9,112,1,2,
/* out0465_em-eta5-phi23*/	4,98,0,6,98,1,3,98,2,15,99,0,2,
/* out0466_em-eta6-phi23*/	4,85,1,1,85,2,10,98,0,9,98,1,1,
/* out0467_em-eta7-phi23*/	3,85,0,9,85,1,7,85,2,3,
/* out0468_em-eta8-phi23*/	3,72,1,5,72,2,8,85,0,2,
/* out0469_em-eta9-phi23*/	2,72,0,5,72,1,8,
/* out0470_em-eta10-phi23*/	8,54,4,1,54,5,13,55,0,2,55,4,2,55,5,12,71,0,1,71,2,1,72,0,1,
/* out0471_em-eta11-phi23*/	4,54,4,11,54,5,3,55,0,12,55,1,8,
/* out0472_em-eta12-phi23*/	6,34,5,2,35,5,2,53,2,12,53,5,1,54,1,4,55,1,8,
/* out0473_em-eta13-phi23*/	4,34,4,5,34,5,12,53,2,3,53,3,4,
/* out0474_em-eta14-phi23*/	4,33,5,3,34,4,11,35,0,1,35,1,5,
/* out0475_em-eta15-phi23*/	3,33,2,9,33,5,5,35,1,3,
/* out0476_em-eta16-phi23*/	3,15,5,1,33,2,6,33,3,6,
/* out0477_em-eta17-phi23*/	3,15,4,5,32,3,1,33,3,6,
/* out0478_em-eta18-phi23*/	3,14,2,8,14,3,2,15,4,3,
/* out0479_em-eta19-phi23*/	5,13,1,10,13,3,10,14,1,5,14,3,9,14,4,1,
/* out0480_em-eta0-phi24*/	0,
/* out0481_em-eta1-phi24*/	0,
/* out0482_em-eta2-phi24*/	1,113,2,1,
/* out0483_em-eta3-phi24*/	6,100,1,4,112,0,11,112,1,2,112,2,14,113,0,9,113,2,2,
/* out0484_em-eta4-phi24*/	5,99,0,2,99,1,12,99,2,10,100,1,3,112,0,5,
/* out0485_em-eta5-phi24*/	5,86,1,10,86,2,1,98,0,1,99,0,12,99,2,2,
/* out0486_em-eta6-phi24*/	4,85,2,2,86,0,13,86,1,6,86,2,1,
/* out0487_em-eta7-phi24*/	4,73,1,8,73,2,3,85,0,5,85,2,1,
/* out0488_em-eta8-phi24*/	3,72,0,1,72,2,8,73,1,6,
/* out0489_em-eta9-phi24*/	2,56,1,3,72,0,9,
/* out0490_em-eta10-phi24*/	5,55,2,16,55,3,8,55,4,9,55,5,4,56,0,1,
/* out0491_em-eta11-phi24*/	7,54,0,3,54,1,3,54,2,16,54,3,5,55,0,2,55,3,1,55,4,5,
/* out0492_em-eta12-phi24*/	4,35,2,5,35,5,8,54,0,6,54,1,9,
/* out0493_em-eta13-phi24*/	4,34,5,2,35,0,7,35,4,10,35,5,6,
/* out0494_em-eta14-phi24*/	4,34,1,2,34,2,6,35,0,8,35,1,4,
/* out0495_em-eta15-phi24*/	4,16,5,3,33,2,1,34,1,8,35,1,4,
/* out0496_em-eta16-phi24*/	3,15,5,10,16,0,1,16,5,4,
/* out0497_em-eta17-phi24*/	3,15,4,4,15,5,5,16,0,3,
/* out0498_em-eta18-phi24*/	2,15,4,4,16,1,6,
/* out0499_em-eta19-phi24*/	5,13,1,2,13,3,2,14,1,1,14,3,4,16,1,4,
/* out0500_em-eta0-phi25*/	0,
/* out0501_em-eta1-phi25*/	0,
/* out0502_em-eta2-phi25*/	3,101,0,3,101,1,3,113,2,7,
/* out0503_em-eta3-phi25*/	6,100,0,3,100,1,3,100,2,16,101,0,10,113,0,7,113,2,6,
/* out0504_em-eta4-phi25*/	5,87,1,10,87,2,1,99,2,3,100,0,12,100,1,6,
/* out0505_em-eta5-phi25*/	6,74,2,1,86,2,5,87,0,13,87,1,6,87,2,1,99,2,1,
/* out0506_em-eta6-phi25*/	5,73,2,1,74,1,9,74,2,1,86,0,3,86,2,9,
/* out0507_em-eta7-phi25*/	4,73,0,4,73,1,1,73,2,12,74,1,1,
/* out0508_em-eta8-phi25*/	3,56,1,4,73,0,10,73,1,1,
/* out0509_em-eta9-phi25*/	3,56,0,3,56,1,9,56,2,1,
/* out0510_em-eta10-phi25*/	4,36,4,3,54,3,1,55,3,7,56,0,8,
/* out0511_em-eta11-phi25*/	4,36,4,9,37,1,11,54,0,4,54,3,10,
/* out0512_em-eta12-phi25*/	5,35,2,10,35,3,1,36,1,10,37,1,4,54,0,3,
/* out0513_em-eta13-phi25*/	5,34,2,3,34,3,3,35,2,1,35,3,12,35,4,6,
/* out0514_em-eta14-phi25*/	4,34,0,5,34,1,3,34,2,7,34,3,5,
/* out0515_em-eta15-phi25*/	4,16,2,5,16,5,3,34,0,6,34,1,3,
/* out0516_em-eta16-phi25*/	4,16,0,1,16,2,1,16,4,6,16,5,6,
/* out0517_em-eta17-phi25*/	3,15,2,2,16,0,8,16,4,3,
/* out0518_em-eta18-phi25*/	4,15,1,2,15,2,2,16,0,3,16,1,3,
/* out0519_em-eta19-phi25*/	2,15,1,5,16,1,3,
/* out0520_em-eta0-phi26*/	0,
/* out0521_em-eta1-phi26*/	0,
/* out0522_em-eta2-phi26*/	2,101,1,10,101,2,1,
/* out0523_em-eta3-phi26*/	7,88,1,9,88,2,4,89,0,7,100,0,1,101,0,3,101,1,3,101,2,15,
/* out0524_em-eta4-phi26*/	5,75,1,2,87,2,6,88,0,14,88,1,7,88,2,3,
/* out0525_em-eta5-phi26*/	5,74,2,4,75,0,4,75,1,8,87,0,3,87,2,8,
/* out0526_em-eta6-phi26*/	3,74,0,8,74,1,4,74,2,10,
/* out0527_em-eta7-phi26*/	5,57,1,4,57,2,6,73,0,1,74,0,5,74,1,2,
/* out0528_em-eta8-phi26*/	3,56,2,2,57,1,12,73,0,1,
/* out0529_em-eta9-phi26*/	2,38,1,1,56,2,11,
/* out0530_em-eta10-phi26*/	6,36,4,2,36,5,11,37,5,4,38,1,1,56,0,4,56,2,2,
/* out0531_em-eta11-phi26*/	7,36,2,2,36,4,2,36,5,5,37,0,16,37,1,1,37,4,7,37,5,2,
/* out0532_em-eta12-phi26*/	4,36,0,8,36,1,6,36,2,12,36,3,3,
/* out0533_em-eta13-phi26*/	5,17,5,5,18,5,4,34,3,5,35,3,3,36,0,7,
/* out0534_em-eta14-phi26*/	4,17,4,7,17,5,7,34,0,4,34,3,3,
/* out0535_em-eta15-phi26*/	3,16,2,8,17,4,8,34,0,1,
/* out0536_em-eta16-phi26*/	3,16,2,2,16,3,8,16,4,4,
/* out0537_em-eta17-phi26*/	3,15,2,8,15,3,1,16,4,3,
/* out0538_em-eta18-phi26*/	3,15,0,2,15,1,4,15,2,4,
/* out0539_em-eta19-phi26*/	2,15,0,1,15,1,5,
/* out0540_em-eta0-phi27*/	0,
/* out0541_em-eta1-phi27*/	0,
/* out0542_em-eta2-phi27*/	0,
/* out0543_em-eta3-phi27*/	4,76,1,7,88,2,3,89,0,9,89,2,16,
/* out0544_em-eta4-phi27*/	6,75,1,3,75,2,4,76,0,8,76,1,9,88,0,2,88,2,6,
/* out0545_em-eta5-phi27*/	4,58,2,1,75,0,11,75,1,3,75,2,12,
/* out0546_em-eta6-phi27*/	4,58,1,10,58,2,7,74,0,3,75,0,1,
/* out0547_em-eta7-phi27*/	3,57,0,2,57,2,10,58,1,6,
/* out0548_em-eta8-phi27*/	2,38,1,1,57,0,13,
/* out0549_em-eta9-phi27*/	2,38,1,12,57,0,1,
/* out0550_em-eta10-phi27*/	4,37,2,1,37,5,5,38,0,8,38,1,1,
/* out0551_em-eta11-phi27*/	4,37,2,15,37,3,7,37,4,7,37,5,5,
/* out0552_em-eta12-phi27*/	5,18,2,3,36,2,2,36,3,13,37,3,9,37,4,2,
/* out0553_em-eta13-phi27*/	5,17,5,1,18,2,5,18,4,5,18,5,12,36,0,1,
/* out0554_em-eta14-phi27*/	3,17,5,3,18,0,14,18,4,3,
/* out0555_em-eta15-phi27*/	3,17,4,1,18,0,2,18,1,13,
/* out0556_em-eta16-phi27*/	3,15,3,4,16,3,8,18,1,3,
/* out0557_em-eta17-phi27*/	2,15,0,1,15,3,11,
/* out0558_em-eta18-phi27*/	1,15,0,10,
/* out0559_em-eta19-phi27*/	1,15,0,2,
/* out0560_em-eta0-phi28*/	0,
/* out0561_em-eta1-phi28*/	0,
/* out0562_em-eta2-phi28*/	0,
/* out0563_em-eta3-phi28*/	1,76,2,7,
/* out0564_em-eta4-phi28*/	2,76,0,8,76,2,9,
/* out0565_em-eta5-phi28*/	1,58,2,1,
/* out0566_em-eta6-phi28*/	2,58,0,10,58,2,7,
/* out0567_em-eta7-phi28*/	1,58,0,6,
/* out0568_em-eta8-phi28*/	1,38,2,1,
/* out0569_em-eta9-phi28*/	1,38,2,12,
/* out0570_em-eta10-phi28*/	2,38,0,8,38,2,1,
/* out0571_em-eta11-phi28*/	0,
/* out0572_em-eta12-phi28*/	1,18,2,3,
/* out0573_em-eta13-phi28*/	4,17,3,1,18,2,5,18,3,12,18,4,5,
/* out0574_em-eta14-phi28*/	3,17,2,14,17,3,3,18,4,3,
/* out0575_em-eta15-phi28*/	3,17,0,1,17,1,13,17,2,2,
/* out0576_em-eta16-phi28*/	1,17,1,3,
/* out0577_em-eta17-phi28*/	0,
/* out0578_em-eta18-phi28*/	0,
/* out0579_em-eta19-phi28*/	0,
/* out0580_em-eta0-phi29*/	0,
/* out0581_em-eta1-phi29*/	0,
/* out0582_em-eta2-phi29*/	0,
/* out0583_em-eta3-phi29*/	0,
/* out0584_em-eta4-phi29*/	0,
/* out0585_em-eta5-phi29*/	0,
/* out0586_em-eta6-phi29*/	0,
/* out0587_em-eta7-phi29*/	0,
/* out0588_em-eta8-phi29*/	0,
/* out0589_em-eta9-phi29*/	1,38,2,1,
/* out0590_em-eta10-phi29*/	1,38,2,1,
/* out0591_em-eta11-phi29*/	0,
/* out0592_em-eta12-phi29*/	0,
/* out0593_em-eta13-phi29*/	2,17,3,5,18,3,4,
/* out0594_em-eta14-phi29*/	2,17,0,7,17,3,7,
/* out0595_em-eta15-phi29*/	1,17,0,8,
/* out0596_em-eta16-phi29*/	0,
/* out0597_em-eta17-phi29*/	0,
/* out0598_em-eta18-phi29*/	0,
/* out0599_em-eta19-phi29*/	0
};