parameter integer matrixH [0:6371] = {
/* num inputs = 251(in0-in250) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1963 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	1,99,0,2,
/* out0002_em-eta2-phi0*/	2,99,0,14,99,1,11,
/* out0003_em-eta3-phi0*/	2,98,0,13,99,1,5,
/* out0004_em-eta4-phi0*/	5,87,2,2,94,0,1,94,1,5,98,0,3,98,1,13,
/* out0005_em-eta5-phi0*/	7,86,0,1,87,2,1,94,0,8,94,1,10,94,2,14,97,0,15,98,1,3,
/* out0006_em-eta6-phi0*/	8,86,0,1,93,0,7,93,1,14,93,2,4,94,0,7,94,2,1,97,0,1,97,1,15,
/* out0007_em-eta7-phi0*/	7,92,0,2,92,1,9,93,0,9,93,2,9,96,0,16,96,1,1,97,1,1,
/* out0008_em-eta8-phi0*/	5,92,0,7,92,1,4,92,2,8,96,1,15,96,2,1,
/* out0009_em-eta9-phi0*/	5,91,0,3,91,1,9,92,0,7,92,2,3,96,2,15,
/* out0010_em-eta10-phi0*/	4,91,0,6,91,1,1,91,2,6,95,0,14,
/* out0011_em-eta11-phi0*/	7,90,0,2,90,1,6,91,0,7,91,2,2,127,2,6,95,0,2,95,1,16,
/* out0012_em-eta12-phi0*/	7,90,0,12,90,1,1,90,2,2,126,0,1,126,1,1,127,1,2,127,2,6,
/* out0013_em-eta13-phi0*/	5,89,0,1,89,1,2,90,0,2,90,2,4,126,0,9,
/* out0014_em-eta14-phi0*/	4,89,0,3,89,1,3,126,0,4,126,2,1,
/* out0015_em-eta15-phi0*/	3,89,0,10,89,2,1,125,0,4,
/* out0016_em-eta16-phi0*/	4,88,0,1,89,0,2,89,2,3,125,0,5,
/* out0017_em-eta17-phi0*/	3,88,0,3,88,1,2,125,0,1,
/* out0018_em-eta18-phi0*/	2,88,0,4,124,0,3,
/* out0019_em-eta19-phi0*/	2,88,0,1,124,0,2,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	1,99,3,2,
/* out0022_em-eta2-phi1*/	2,99,2,11,99,3,14,
/* out0023_em-eta3-phi1*/	2,98,3,13,99,2,5,
/* out0024_em-eta4-phi1*/	4,87,1,5,87,2,9,98,2,13,98,3,3,
/* out0025_em-eta5-phi1*/	9,86,0,7,86,1,12,86,2,1,87,1,9,87,2,4,94,1,1,94,2,1,97,3,15,98,2,3,
/* out0026_em-eta6-phi1*/	8,85,0,1,85,1,5,86,0,7,86,2,9,93,1,2,93,2,2,97,2,15,97,3,1,
/* out0027_em-eta7-phi1*/	8,85,0,14,85,1,2,85,2,3,92,1,1,93,2,1,96,4,1,96,5,16,97,2,1,
/* out0028_em-eta8-phi1*/	8,84,0,6,84,1,3,85,0,1,85,2,2,92,1,2,92,2,5,96,3,1,96,4,15,
/* out0029_em-eta9-phi1*/	4,84,0,9,84,2,1,91,1,5,96,3,15,
/* out0030_em-eta10-phi1*/	4,83,0,4,91,1,1,91,2,7,95,3,14,
/* out0031_em-eta11-phi1*/	7,83,0,4,90,1,6,91,2,1,127,1,4,127,2,4,95,2,16,95,3,2,
/* out0032_em-eta12-phi1*/	5,90,1,3,90,2,6,122,0,1,126,1,5,127,1,9,
/* out0033_em-eta13-phi1*/	6,82,0,2,89,1,2,90,2,4,126,0,2,126,1,7,126,2,3,
/* out0034_em-eta14-phi1*/	3,89,1,6,125,1,2,126,2,7,
/* out0035_em-eta15-phi1*/	4,89,1,1,89,2,4,125,0,2,125,1,7,
/* out0036_em-eta16-phi1*/	4,88,1,1,89,2,4,125,0,3,125,2,3,
/* out0037_em-eta17-phi1*/	5,88,0,1,88,1,5,124,1,2,125,0,1,125,2,3,
/* out0038_em-eta18-phi1*/	4,88,0,3,88,1,1,124,0,5,124,1,1,
/* out0039_em-eta19-phi1*/	1,124,0,2,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	1,104,0,2,
/* out0042_em-eta2-phi2*/	2,104,0,14,104,1,11,
/* out0043_em-eta3-phi2*/	2,103,0,13,104,1,5,
/* out0044_em-eta4-phi2*/	5,80,0,11,80,2,4,87,1,2,103,0,3,103,1,13,
/* out0045_em-eta5-phi2*/	8,79,1,4,80,0,3,80,1,10,80,2,12,86,1,4,86,2,1,102,0,15,103,1,3,
/* out0046_em-eta6-phi2*/	7,79,0,15,79,1,2,79,2,1,85,1,4,86,2,5,102,0,1,102,1,15,
/* out0047_em-eta7-phi2*/	9,78,0,5,78,1,1,79,0,1,79,2,1,85,1,5,85,2,10,101,0,16,101,1,1,102,1,1,
/* out0048_em-eta8-phi2*/	6,78,0,3,84,1,13,84,2,1,85,2,1,101,1,15,101,2,1,
/* out0049_em-eta9-phi2*/	4,83,1,1,84,0,1,84,2,13,101,2,15,
/* out0050_em-eta10-phi2*/	4,83,0,3,83,1,10,83,2,1,100,0,14,
/* out0051_em-eta11-phi2*/	7,83,0,5,83,2,6,122,0,3,122,1,6,127,1,1,100,0,2,100,1,16,
/* out0052_em-eta12-phi2*/	6,82,0,3,82,1,4,83,2,1,122,0,11,122,1,1,122,2,2,
/* out0053_em-eta13-phi2*/	7,82,0,7,121,0,2,121,1,1,122,0,1,122,2,1,126,1,3,126,2,3,
/* out0054_em-eta14-phi2*/	6,82,0,3,82,2,1,89,1,2,121,0,7,125,1,1,126,2,2,
/* out0055_em-eta15-phi2*/	5,81,0,2,89,2,3,121,0,1,125,1,6,125,2,1,
/* out0056_em-eta16-phi2*/	3,81,0,3,89,2,1,125,2,7,
/* out0057_em-eta17-phi2*/	5,81,0,1,88,1,4,120,0,1,124,1,4,125,2,2,
/* out0058_em-eta18-phi2*/	4,88,0,2,88,1,2,124,0,2,124,1,4,
/* out0059_em-eta19-phi2*/	1,124,0,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	1,104,3,2,
/* out0062_em-eta2-phi3*/	2,104,2,11,104,3,14,
/* out0063_em-eta3-phi3*/	2,103,3,13,104,2,5,
/* out0064_em-eta4-phi3*/	4,74,1,3,80,0,2,103,2,13,103,3,3,
/* out0065_em-eta5-phi3*/	7,74,0,15,74,1,4,74,2,2,79,1,4,80,1,6,102,3,15,103,2,3,
/* out0066_em-eta6-phi3*/	7,73,0,5,74,0,1,74,2,1,79,1,6,79,2,13,102,2,15,102,3,1,
/* out0067_em-eta7-phi3*/	8,73,0,1,78,0,4,78,1,14,78,2,3,79,2,1,101,4,1,101,5,16,102,2,1,
/* out0068_em-eta8-phi3*/	6,77,0,1,77,1,4,78,0,4,78,2,8,101,3,1,101,4,15,
/* out0069_em-eta9-phi3*/	4,77,0,12,77,1,2,84,2,1,101,3,15,
/* out0070_em-eta10-phi3*/	6,76,0,1,77,0,3,77,2,1,83,1,5,83,2,2,100,3,14,
/* out0071_em-eta11-phi3*/	5,76,0,4,83,2,6,122,1,7,100,2,16,100,3,2,
/* out0072_em-eta12-phi3*/	4,82,1,8,122,1,2,122,2,11,123,1,1,
/* out0073_em-eta13-phi3*/	5,82,0,1,82,1,2,82,2,5,121,1,9,122,2,2,
/* out0074_em-eta14-phi3*/	5,81,1,2,82,2,4,121,0,4,121,1,2,121,2,3,
/* out0075_em-eta15-phi3*/	5,81,0,2,81,1,3,120,1,2,121,0,2,121,2,4,
/* out0076_em-eta16-phi3*/	3,81,0,4,120,0,5,120,1,1,
/* out0077_em-eta17-phi3*/	3,81,0,3,120,0,5,124,1,1,
/* out0078_em-eta18-phi3*/	5,88,0,1,88,1,1,120,0,1,124,0,1,124,1,4,
/* out0079_em-eta19-phi3*/	0,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	1,109,0,2,
/* out0082_em-eta2-phi4*/	2,109,0,14,109,1,11,
/* out0083_em-eta3-phi4*/	2,108,0,13,109,1,5,
/* out0084_em-eta4-phi4*/	3,74,1,3,108,0,3,108,1,13,
/* out0085_em-eta5-phi4*/	7,73,1,1,74,1,6,74,2,13,75,1,9,75,2,2,107,0,15,108,1,3,
/* out0086_em-eta6-phi4*/	5,73,0,6,73,1,14,73,2,6,107,0,1,107,1,15,
/* out0087_em-eta7-phi4*/	9,72,0,3,72,1,5,73,0,4,73,2,6,78,1,1,78,2,3,106,0,16,106,1,1,107,1,1,
/* out0088_em-eta8-phi4*/	5,72,0,11,77,1,5,78,2,2,106,1,15,106,2,1,
/* out0089_em-eta9-phi4*/	3,77,1,5,77,2,10,106,2,15,
/* out0090_em-eta10-phi4*/	3,76,1,8,77,2,5,105,0,14,
/* out0091_em-eta11-phi4*/	6,76,0,7,76,1,2,76,2,1,123,2,4,105,0,2,105,1,16,
/* out0092_em-eta12-phi4*/	7,76,0,4,76,2,2,82,1,2,82,2,1,123,0,1,123,1,9,123,2,4,
/* out0093_em-eta13-phi4*/	5,60,1,3,82,2,4,121,1,4,123,0,1,123,1,6,
/* out0094_em-eta14-phi4*/	5,60,1,2,81,1,3,82,2,1,116,0,2,121,2,7,
/* out0095_em-eta15-phi4*/	4,81,1,5,116,0,1,120,1,5,121,2,2,
/* out0096_em-eta16-phi4*/	5,81,0,1,81,2,4,120,0,1,120,1,5,120,2,1,
/* out0097_em-eta17-phi4*/	3,81,2,4,120,0,2,120,2,3,
/* out0098_em-eta18-phi4*/	2,120,0,1,120,2,2,
/* out0099_em-eta19-phi4*/	0,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	1,109,3,2,
/* out0102_em-eta2-phi5*/	2,109,2,11,109,3,14,
/* out0103_em-eta3-phi5*/	2,108,3,13,109,2,5,
/* out0104_em-eta4-phi5*/	3,75,2,2,108,2,13,108,3,3,
/* out0105_em-eta5-phi5*/	5,75,0,13,75,1,5,75,2,12,107,3,15,108,2,3,
/* out0106_em-eta6-phi5*/	8,68,0,9,68,1,8,73,1,1,73,2,3,75,0,3,75,1,2,107,2,15,107,3,1,
/* out0107_em-eta7-phi5*/	7,68,0,7,72,1,11,72,2,2,73,2,1,106,4,1,106,5,16,107,2,1,
/* out0108_em-eta8-phi5*/	5,66,2,2,72,0,2,72,2,14,106,3,1,106,4,15,
/* out0109_em-eta9-phi5*/	3,66,1,9,66,2,5,106,3,15,
/* out0110_em-eta10-phi5*/	3,66,1,7,76,1,5,105,3,14,
/* out0111_em-eta11-phi5*/	5,76,1,1,76,2,9,123,2,3,105,2,16,105,3,2,
/* out0112_em-eta12-phi5*/	4,60,2,5,76,2,4,123,0,8,123,2,5,
/* out0113_em-eta13-phi5*/	4,60,1,5,60,2,2,116,1,5,123,0,6,
/* out0114_em-eta14-phi5*/	3,60,1,6,116,0,7,116,1,3,
/* out0115_em-eta15-phi5*/	4,81,1,3,81,2,2,116,0,6,120,1,1,
/* out0116_em-eta16-phi5*/	3,81,2,4,120,1,2,120,2,4,
/* out0117_em-eta17-phi5*/	2,81,2,2,120,2,5,
/* out0118_em-eta18-phi5*/	1,120,2,1,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	1,114,0,2,
/* out0122_em-eta2-phi6*/	2,114,0,14,114,1,11,
/* out0123_em-eta3-phi6*/	2,113,0,13,114,1,5,
/* out0124_em-eta4-phi6*/	3,70,1,2,113,0,3,113,1,13,
/* out0125_em-eta5-phi6*/	5,70,0,13,70,1,12,70,2,5,112,0,15,113,1,3,
/* out0126_em-eta6-phi6*/	8,68,1,8,68,2,9,69,1,3,69,2,1,70,0,3,70,2,2,112,0,1,112,1,15,
/* out0127_em-eta7-phi6*/	7,67,1,3,67,2,11,68,2,7,69,1,1,111,0,16,111,1,1,112,1,1,
/* out0128_em-eta8-phi6*/	5,66,2,3,67,0,2,67,1,13,111,1,15,111,2,1,
/* out0129_em-eta9-phi6*/	3,66,0,9,66,2,6,111,2,15,
/* out0130_em-eta10-phi6*/	3,61,2,5,66,0,7,110,0,14,
/* out0131_em-eta11-phi6*/	5,61,1,9,61,2,1,118,1,3,110,0,2,110,1,16,
/* out0132_em-eta12-phi6*/	4,60,2,5,61,1,4,118,0,8,118,1,5,
/* out0133_em-eta13-phi6*/	4,60,0,4,60,2,3,116,1,5,118,0,6,
/* out0134_em-eta14-phi6*/	3,60,0,6,116,1,3,116,2,6,
/* out0135_em-eta15-phi6*/	5,53,1,2,53,2,3,60,0,1,115,2,1,116,2,6,
/* out0136_em-eta16-phi6*/	3,53,1,4,115,1,4,115,2,2,
/* out0137_em-eta17-phi6*/	2,53,1,2,115,1,5,
/* out0138_em-eta18-phi6*/	1,115,1,1,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	1,114,3,2,
/* out0142_em-eta2-phi7*/	2,114,2,11,114,3,14,
/* out0143_em-eta3-phi7*/	2,113,3,13,114,2,5,
/* out0144_em-eta4-phi7*/	3,71,2,3,113,2,13,113,3,3,
/* out0145_em-eta5-phi7*/	7,69,2,1,70,1,2,70,2,9,71,1,13,71,2,6,112,3,15,113,2,3,
/* out0146_em-eta6-phi7*/	5,69,0,6,69,1,6,69,2,14,112,2,15,112,3,1,
/* out0147_em-eta7-phi7*/	9,63,1,3,63,2,1,67,0,3,67,2,5,69,0,4,69,1,6,111,4,1,111,5,16,112,2,1,
/* out0148_em-eta8-phi7*/	5,62,2,5,63,1,2,67,0,11,111,3,1,111,4,15,
/* out0149_em-eta9-phi7*/	3,62,1,10,62,2,5,111,3,15,
/* out0150_em-eta10-phi7*/	3,61,2,8,62,1,5,110,3,14,
/* out0151_em-eta11-phi7*/	6,61,0,7,61,1,1,61,2,2,118,1,4,110,2,16,110,3,2,
/* out0152_em-eta12-phi7*/	8,54,1,1,54,2,2,60,2,1,61,0,4,61,1,2,118,0,1,118,1,4,118,2,9,
/* out0153_em-eta13-phi7*/	5,54,1,4,60,0,3,117,2,4,118,0,1,118,2,6,
/* out0154_em-eta14-phi7*/	5,53,2,3,54,1,1,60,0,2,116,2,3,117,1,7,
/* out0155_em-eta15-phi7*/	4,53,2,5,115,2,5,116,2,1,117,1,2,
/* out0156_em-eta16-phi7*/	5,53,0,1,53,1,4,115,0,1,115,1,1,115,2,5,
/* out0157_em-eta17-phi7*/	3,53,1,4,115,0,2,115,1,3,
/* out0158_em-eta18-phi7*/	2,115,0,1,115,1,2,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	1,119,0,2,
/* out0162_em-eta2-phi8*/	2,119,0,14,119,1,11,
/* out0163_em-eta3-phi8*/	2,118,0,13,119,1,5,
/* out0164_em-eta4-phi8*/	4,65,0,2,71,2,3,118,0,3,118,1,13,
/* out0165_em-eta5-phi8*/	8,64,2,4,65,0,1,65,2,7,71,0,15,71,1,2,71,2,4,117,0,15,118,1,3,
/* out0166_em-eta6-phi8*/	7,64,1,13,64,2,6,69,0,5,71,0,1,71,1,1,117,0,1,117,1,15,
/* out0167_em-eta7-phi8*/	8,63,0,4,63,1,3,63,2,14,64,1,1,69,0,1,116,0,16,116,1,1,117,1,1,
/* out0168_em-eta8-phi8*/	6,62,0,1,62,2,4,63,0,4,63,1,8,116,1,15,116,2,1,
/* out0169_em-eta9-phi8*/	4,56,1,1,62,0,12,62,2,2,116,2,15,
/* out0170_em-eta10-phi8*/	6,55,1,2,55,2,5,61,0,1,62,0,3,62,1,1,115,0,14,
/* out0171_em-eta11-phi8*/	5,55,1,6,61,0,4,119,2,7,115,0,2,115,1,16,
/* out0172_em-eta12-phi8*/	4,54,2,8,118,2,1,119,1,11,119,2,2,
/* out0173_em-eta13-phi8*/	5,54,0,1,54,1,5,54,2,2,117,2,9,119,1,2,
/* out0174_em-eta14-phi8*/	5,53,2,2,54,1,4,117,0,4,117,1,3,117,2,2,
/* out0175_em-eta15-phi8*/	5,53,0,2,53,2,3,115,2,2,117,0,2,117,1,4,
/* out0176_em-eta16-phi8*/	3,53,0,4,115,0,5,115,2,1,
/* out0177_em-eta17-phi8*/	2,53,0,3,115,0,5,
/* out0178_em-eta18-phi8*/	3,46,1,2,111,1,5,115,0,1,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	1,119,3,2,
/* out0182_em-eta2-phi9*/	2,119,2,11,119,3,14,
/* out0183_em-eta3-phi9*/	2,118,3,13,119,2,5,
/* out0184_em-eta4-phi9*/	5,59,1,2,65,0,9,65,1,4,118,2,13,118,3,3,
/* out0185_em-eta5-phi9*/	8,58,1,1,58,2,4,64,2,4,65,0,4,65,1,12,65,2,9,117,3,15,118,2,3,
/* out0186_em-eta6-phi9*/	7,57,2,4,58,1,5,64,0,15,64,1,1,64,2,2,117,2,15,117,3,1,
/* out0187_em-eta7-phi9*/	9,57,1,10,57,2,5,63,0,5,63,2,1,64,0,1,64,1,1,116,4,1,116,5,16,117,2,1,
/* out0188_em-eta8-phi9*/	6,56,1,1,56,2,13,57,1,1,63,0,3,116,3,1,116,4,15,
/* out0189_em-eta9-phi9*/	4,55,2,1,56,0,1,56,1,13,116,3,15,
/* out0190_em-eta10-phi9*/	4,55,0,3,55,1,1,55,2,10,115,3,14,
/* out0191_em-eta11-phi9*/	7,55,0,5,55,1,6,114,1,1,119,0,3,119,2,6,115,2,16,115,3,2,
/* out0192_em-eta12-phi9*/	6,54,0,3,54,2,4,55,1,1,119,0,11,119,1,2,119,2,1,
/* out0193_em-eta13-phi9*/	7,54,0,7,113,1,3,113,2,3,117,0,2,117,2,1,119,0,1,119,1,1,
/* out0194_em-eta14-phi9*/	6,47,2,2,54,0,3,54,1,1,112,2,1,113,1,2,117,0,7,
/* out0195_em-eta15-phi9*/	5,47,1,3,53,0,2,112,1,1,112,2,6,117,0,1,
/* out0196_em-eta16-phi9*/	3,47,1,1,53,0,3,112,1,7,
/* out0197_em-eta17-phi9*/	6,46,1,4,53,0,1,111,1,1,111,2,2,112,1,2,115,0,1,
/* out0198_em-eta18-phi9*/	3,46,1,3,111,1,5,111,2,1,
/* out0199_em-eta19-phi9*/	1,111,1,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	1,124,0,2,
/* out0202_em-eta2-phi10*/	2,124,0,14,124,1,11,
/* out0203_em-eta3-phi10*/	2,123,0,13,124,1,5,
/* out0204_em-eta4-phi10*/	4,59,0,9,59,1,5,123,0,3,123,1,13,
/* out0205_em-eta5-phi10*/	9,52,1,1,52,2,1,58,0,7,58,1,1,58,2,12,59,0,4,59,1,9,122,0,15,123,1,3,
/* out0206_em-eta6-phi10*/	8,51,1,2,51,2,2,57,0,1,57,2,5,58,0,7,58,1,9,122,0,1,122,1,15,
/* out0207_em-eta7-phi10*/	8,50,2,1,51,1,1,57,0,14,57,1,3,57,2,2,121,0,16,121,1,1,122,1,1,
/* out0208_em-eta8-phi10*/	8,50,1,5,50,2,2,56,0,6,56,2,3,57,0,1,57,1,2,121,1,15,121,2,1,
/* out0209_em-eta9-phi10*/	4,49,2,5,56,0,9,56,1,1,121,2,15,
/* out0210_em-eta10-phi10*/	4,49,1,7,49,2,1,55,0,4,120,0,14,
/* out0211_em-eta11-phi10*/	7,48,2,6,49,1,1,55,0,4,114,0,4,114,1,4,120,0,2,120,1,16,
/* out0212_em-eta12-phi10*/	5,48,1,6,48,2,3,113,2,5,114,1,9,119,0,1,
/* out0213_em-eta13-phi10*/	6,47,2,2,48,1,4,54,0,2,113,0,2,113,1,3,113,2,7,
/* out0214_em-eta14-phi10*/	3,47,2,6,112,2,2,113,1,7,
/* out0215_em-eta15-phi10*/	4,47,1,4,47,2,1,112,0,2,112,2,7,
/* out0216_em-eta16-phi10*/	4,46,2,1,47,1,4,112,0,3,112,1,3,
/* out0217_em-eta17-phi10*/	5,46,1,1,46,2,4,111,2,3,112,0,1,112,1,3,
/* out0218_em-eta18-phi10*/	3,46,1,3,111,1,1,111,2,6,
/* out0219_em-eta19-phi10*/	1,111,1,2,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	1,124,3,2,
/* out0222_em-eta2-phi11*/	2,124,2,11,124,3,14,
/* out0223_em-eta3-phi11*/	2,123,3,13,124,2,5,
/* out0224_em-eta4-phi11*/	5,52,0,1,52,2,5,59,0,2,123,2,13,123,3,3,
/* out0225_em-eta5-phi11*/	7,52,0,8,52,1,14,52,2,10,58,0,1,59,0,1,122,3,15,123,2,3,
/* out0226_em-eta6-phi11*/	7,51,0,6,51,1,4,51,2,14,52,1,1,58,0,1,122,2,15,122,3,1,
/* out0227_em-eta7-phi11*/	7,50,0,2,50,2,9,51,0,2,51,1,9,121,4,1,121,5,16,122,2,1,
/* out0228_em-eta8-phi11*/	5,50,0,7,50,1,8,50,2,4,121,3,1,121,4,15,
/* out0229_em-eta9-phi11*/	4,49,0,3,49,2,9,50,1,3,121,3,15,
/* out0230_em-eta10-phi11*/	4,49,0,5,49,1,6,49,2,1,120,3,14,
/* out0231_em-eta11-phi11*/	6,48,0,2,48,2,6,49,1,2,114,0,6,120,2,16,120,3,2,
/* out0232_em-eta12-phi11*/	8,48,0,5,48,1,2,48,2,1,110,0,6,113,0,1,113,2,1,114,0,6,114,1,2,
/* out0233_em-eta13-phi11*/	5,47,2,2,48,0,1,48,1,4,110,0,2,113,0,9,
/* out0234_em-eta14-phi11*/	5,47,0,3,47,2,3,109,0,4,113,0,4,113,1,1,
/* out0235_em-eta15-phi11*/	4,47,0,4,47,1,1,109,0,3,112,0,4,
/* out0236_em-eta16-phi11*/	4,47,0,1,47,1,3,108,0,1,112,0,5,
/* out0237_em-eta17-phi11*/	3,46,2,5,108,0,4,112,0,1,
/* out0238_em-eta18-phi11*/	4,46,1,2,46,2,2,108,0,3,111,2,3,
/* out0239_em-eta19-phi11*/	2,111,1,1,111,2,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	1,129,0,2,
/* out0242_em-eta2-phi12*/	2,129,0,14,129,1,11,
/* out0243_em-eta3-phi12*/	2,128,0,13,129,1,5,
/* out0244_em-eta4-phi12*/	4,45,0,9,45,2,1,128,0,3,128,1,13,
/* out0245_em-eta5-phi12*/	7,44,0,7,44,1,8,45,0,6,45,2,8,52,0,7,127,0,15,128,1,3,
/* out0246_em-eta6-phi12*/	7,43,0,1,43,1,3,44,0,9,44,2,7,51,0,6,127,0,1,127,1,15,
/* out0247_em-eta7-phi12*/	8,43,0,14,43,1,3,43,2,2,50,0,1,51,0,2,126,0,16,126,1,1,127,1,1,
/* out0248_em-eta8-phi12*/	7,42,0,5,42,1,3,43,0,1,43,2,2,50,0,6,126,1,15,126,2,1,
/* out0249_em-eta9-phi12*/	4,42,0,11,42,2,1,49,0,3,126,2,15,
/* out0250_em-eta10-phi12*/	5,41,0,5,41,1,1,42,2,1,49,0,5,125,0,14,
/* out0251_em-eta11-phi12*/	5,41,0,8,48,0,2,110,1,5,125,0,2,125,1,16,
/* out0252_em-eta12-phi12*/	7,40,0,2,41,0,1,41,2,1,48,0,5,110,0,6,110,1,5,110,2,2,
/* out0253_em-eta13-phi12*/	5,40,0,6,48,0,1,109,1,3,110,0,2,110,2,6,
/* out0254_em-eta14-phi12*/	4,40,0,3,47,0,3,109,0,5,109,1,4,
/* out0255_em-eta15-phi12*/	4,39,0,1,47,0,4,109,0,4,109,2,5,
/* out0256_em-eta16-phi12*/	5,39,0,3,47,0,1,108,0,1,108,1,4,109,2,1,
/* out0257_em-eta17-phi12*/	4,39,0,3,46,2,1,108,0,4,108,1,1,
/* out0258_em-eta18-phi12*/	4,46,1,1,46,2,3,108,0,3,108,2,2,
/* out0259_em-eta19-phi12*/	1,108,2,2,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	1,129,3,2,
/* out0262_em-eta2-phi13*/	2,129,2,11,129,3,14,
/* out0263_em-eta3-phi13*/	2,128,3,13,129,2,5,
/* out0264_em-eta4-phi13*/	6,38,0,2,38,1,5,45,0,1,45,2,3,128,2,13,128,3,3,
/* out0265_em-eta5-phi13*/	8,37,1,1,38,0,14,38,1,2,38,2,4,44,1,8,45,2,4,127,3,15,128,2,3,
/* out0266_em-eta6-phi13*/	6,37,0,12,37,1,2,43,1,3,44,2,9,127,2,15,127,3,1,
/* out0267_em-eta7-phi13*/	8,36,0,3,37,0,2,37,2,1,43,1,7,43,2,9,126,4,1,126,5,16,127,2,1,
/* out0268_em-eta8-phi13*/	5,36,0,5,42,1,11,43,2,3,126,3,1,126,4,15,
/* out0269_em-eta9-phi13*/	4,35,0,1,42,1,2,42,2,12,126,3,15,
/* out0270_em-eta10-phi13*/	3,41,1,11,42,2,1,125,3,14,
/* out0271_em-eta11-phi13*/	7,41,0,2,41,1,1,41,2,8,107,0,7,110,1,1,125,2,16,125,3,2,
/* out0272_em-eta12-phi13*/	6,40,1,6,41,2,3,105,0,2,107,0,4,110,1,5,110,2,4,
/* out0273_em-eta13-phi13*/	6,40,0,3,40,1,3,40,2,1,105,0,6,109,1,2,110,2,4,
/* out0274_em-eta14-phi13*/	5,40,0,2,40,2,4,105,0,1,109,1,7,109,2,2,
/* out0275_em-eta15-phi13*/	5,39,0,1,39,1,3,40,2,1,103,0,1,109,2,7,
/* out0276_em-eta16-phi13*/	5,39,0,4,39,1,1,103,0,1,108,1,5,109,2,1,
/* out0277_em-eta17-phi13*/	3,39,0,3,108,1,4,108,2,2,
/* out0278_em-eta18-phi13*/	3,39,0,1,39,2,1,108,2,5,
/* out0279_em-eta19-phi13*/	1,108,2,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	1,134,0,2,
/* out0282_em-eta2-phi14*/	2,134,0,14,134,1,11,
/* out0283_em-eta3-phi14*/	2,133,0,13,134,1,5,
/* out0284_em-eta4-phi14*/	3,38,1,5,133,0,3,133,1,13,
/* out0285_em-eta5-phi14*/	7,32,0,11,32,1,2,37,1,2,38,1,4,38,2,12,132,0,15,133,1,3,
/* out0286_em-eta6-phi14*/	7,31,0,1,32,0,2,37,0,2,37,1,11,37,2,10,132,0,1,132,1,15,
/* out0287_em-eta7-phi14*/	7,31,0,2,36,0,2,36,1,13,37,2,5,131,0,16,131,1,1,132,1,1,
/* out0288_em-eta8-phi14*/	5,35,1,1,36,0,6,36,2,10,131,1,15,131,2,1,
/* out0289_em-eta9-phi14*/	4,35,0,8,35,1,6,42,2,1,131,2,15,
/* out0290_em-eta10-phi14*/	4,35,0,7,35,2,3,41,1,3,130,0,14,
/* out0291_em-eta11-phi14*/	7,34,0,5,34,1,1,41,2,4,107,0,5,107,2,7,130,0,2,130,1,16,
/* out0292_em-eta12-phi14*/	4,34,0,5,40,1,3,105,1,8,107,2,7,
/* out0293_em-eta13-phi14*/	5,40,1,4,40,2,4,105,0,5,105,1,3,105,2,3,
/* out0294_em-eta14-phi14*/	5,33,0,1,40,2,5,103,1,3,105,0,2,105,2,4,
/* out0295_em-eta15-phi14*/	3,39,1,5,103,0,7,103,1,1,
/* out0296_em-eta16-phi14*/	3,39,1,3,39,2,1,103,0,6,
/* out0297_em-eta17-phi14*/	6,39,2,4,102,1,1,103,0,1,103,2,1,108,1,2,108,2,2,
/* out0298_em-eta18-phi14*/	3,39,2,2,102,1,2,108,2,2,
/* out0299_em-eta19-phi14*/	2,102,0,1,102,1,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	1,134,3,2,
/* out0302_em-eta2-phi15*/	2,134,2,11,134,3,14,
/* out0303_em-eta3-phi15*/	2,133,3,13,134,2,5,
/* out0304_em-eta4-phi15*/	4,28,0,10,28,2,3,133,2,13,133,3,3,
/* out0305_em-eta5-phi15*/	8,26,0,2,28,1,1,28,2,13,32,0,2,32,1,14,32,2,10,132,3,15,133,2,3,
/* out0306_em-eta6-phi15*/	8,26,0,1,31,0,5,31,1,13,31,2,1,32,0,1,32,2,6,132,2,15,132,3,1,
/* out0307_em-eta7-phi15*/	8,30,1,3,31,0,8,31,2,7,36,1,3,36,2,1,131,4,1,131,5,16,132,2,1,
/* out0308_em-eta8-phi15*/	6,30,0,11,30,1,1,35,1,1,36,2,5,131,3,1,131,4,15,
/* out0309_em-eta9-phi15*/	4,30,0,2,35,1,8,35,2,5,131,3,15,
/* out0310_em-eta10-phi15*/	4,29,0,1,34,1,3,35,2,8,130,3,14,
/* out0311_em-eta11-phi15*/	8,34,0,2,34,1,8,34,2,1,106,0,8,106,2,6,107,2,2,130,2,16,130,3,2,
/* out0312_em-eta12-phi15*/	5,34,0,4,34,2,5,105,1,3,106,1,2,106,2,10,
/* out0313_em-eta13-phi15*/	7,33,0,2,33,1,3,34,2,1,40,2,1,104,1,3,105,1,2,105,2,6,
/* out0314_em-eta14-phi15*/	4,33,0,6,103,1,5,104,1,2,105,2,3,
/* out0315_em-eta15-phi15*/	4,33,0,3,39,1,2,103,1,5,103,2,2,
/* out0316_em-eta16-phi15*/	3,39,1,2,39,2,2,103,2,6,
/* out0317_em-eta17-phi15*/	3,39,2,4,102,1,4,103,2,1,
/* out0318_em-eta18-phi15*/	3,39,2,1,102,0,1,102,1,4,
/* out0319_em-eta19-phi15*/	1,102,0,4,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	1,139,0,2,
/* out0322_em-eta2-phi16*/	2,139,0,14,139,1,11,
/* out0323_em-eta3-phi16*/	2,138,0,13,139,1,5,
/* out0324_em-eta4-phi16*/	6,27,1,5,27,2,1,28,0,6,28,1,5,138,0,3,138,1,13,
/* out0325_em-eta5-phi16*/	8,26,0,6,26,1,14,26,2,3,27,0,2,27,1,8,28,1,10,137,0,15,138,1,3,
/* out0326_em-eta6-phi16*/	8,25,0,2,25,1,4,26,0,7,26,2,7,31,1,3,31,2,3,137,0,1,137,1,15,
/* out0327_em-eta7-phi16*/	6,25,0,11,30,1,6,31,2,5,136,0,16,136,1,1,137,1,1,
/* out0328_em-eta8-phi16*/	5,30,0,2,30,1,6,30,2,10,136,1,15,136,2,1,
/* out0329_em-eta9-phi16*/	5,29,0,3,29,1,8,30,0,1,30,2,4,136,2,15,
/* out0330_em-eta10-phi16*/	3,29,0,11,29,2,1,135,0,14,
/* out0331_em-eta11-phi16*/	9,14,1,1,29,0,1,29,2,1,34,1,4,34,2,3,106,0,8,106,1,4,135,0,2,135,1,16,
/* out0332_em-eta12-phi16*/	5,14,1,2,33,1,1,34,2,6,104,2,2,106,1,10,
/* out0333_em-eta13-phi16*/	3,33,1,7,104,1,4,104,2,7,
/* out0334_em-eta14-phi16*/	5,33,0,2,33,1,1,33,2,3,104,0,2,104,1,7,
/* out0335_em-eta15-phi16*/	6,33,0,2,33,2,3,98,1,1,103,1,2,103,2,3,104,0,1,
/* out0336_em-eta16-phi16*/	4,0,1,3,39,2,1,98,1,3,103,2,3,
/* out0337_em-eta17-phi16*/	3,0,1,3,102,1,2,102,2,3,
/* out0338_em-eta18-phi16*/	5,0,0,2,0,1,1,102,0,2,102,1,2,102,2,2,
/* out0339_em-eta19-phi16*/	1,102,0,6,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	1,139,3,2,
/* out0342_em-eta2-phi17*/	2,139,2,11,139,3,14,
/* out0343_em-eta3-phi17*/	2,138,3,13,139,2,5,
/* out0344_em-eta4-phi17*/	3,27,2,7,138,2,13,138,3,3,
/* out0345_em-eta5-phi17*/	9,23,0,5,23,1,8,26,1,2,26,2,3,27,0,14,27,1,3,27,2,8,137,3,15,138,2,3,
/* out0346_em-eta6-phi17*/	6,23,0,11,25,1,11,25,2,1,26,2,3,137,2,15,137,3,1,
/* out0347_em-eta7-phi17*/	7,19,2,2,25,0,3,25,1,1,25,2,15,136,4,1,136,5,16,137,2,1,
/* out0348_em-eta8-phi17*/	5,19,1,10,19,2,5,30,2,2,136,3,1,136,4,15,
/* out0349_em-eta9-phi17*/	4,19,1,6,29,1,8,29,2,2,136,3,15,
/* out0350_em-eta10-phi17*/	2,29,2,11,135,3,14,
/* out0351_em-eta11-phi17*/	7,14,1,2,14,2,7,29,2,1,101,0,8,101,2,2,135,2,16,135,3,2,
/* out0352_em-eta12-phi17*/	5,14,1,9,101,0,1,101,1,1,101,2,13,104,2,1,
/* out0353_em-eta13-phi17*/	6,14,1,2,33,1,4,33,2,1,101,2,1,104,0,5,104,2,6,
/* out0354_em-eta14-phi17*/	3,33,2,6,98,2,1,104,0,8,
/* out0355_em-eta15-phi17*/	4,0,1,2,33,2,3,98,1,2,98,2,6,
/* out0356_em-eta16-phi17*/	2,0,1,4,98,1,7,
/* out0357_em-eta17-phi17*/	4,0,0,2,0,1,2,98,1,3,102,2,3,
/* out0358_em-eta18-phi17*/	2,0,0,3,102,2,6,
/* out0359_em-eta19-phi17*/	2,102,0,2,102,2,2,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	1,144,0,2,
/* out0362_em-eta2-phi18*/	2,144,0,14,144,1,11,
/* out0363_em-eta3-phi18*/	2,143,0,13,144,1,5,
/* out0364_em-eta4-phi18*/	3,24,0,8,143,0,3,143,1,13,
/* out0365_em-eta5-phi18*/	9,21,1,3,21,2,2,23,1,8,23,2,5,24,0,7,24,1,9,24,2,16,142,0,15,143,1,3,
/* out0366_em-eta6-phi18*/	6,20,1,1,20,2,11,21,1,3,23,2,11,142,0,1,142,1,15,
/* out0367_em-eta7-phi18*/	7,19,2,3,20,0,3,20,1,15,20,2,1,141,0,16,141,1,1,142,1,1,
/* out0368_em-eta8-phi18*/	5,16,1,2,19,0,10,19,2,6,141,1,15,141,2,1,
/* out0369_em-eta9-phi18*/	4,15,1,2,15,2,8,19,0,6,141,2,15,
/* out0370_em-eta10-phi18*/	3,14,2,1,15,1,11,140,0,14,
/* out0371_em-eta11-phi18*/	7,14,0,2,14,2,8,15,1,1,101,0,7,101,1,3,140,0,2,140,1,16,
/* out0372_em-eta12-phi18*/	3,14,0,8,99,2,1,101,1,11,
/* out0373_em-eta13-phi18*/	6,1,1,1,1,2,4,14,0,3,99,1,5,99,2,6,101,1,1,
/* out0374_em-eta14-phi18*/	3,1,1,6,98,2,1,99,1,8,
/* out0375_em-eta15-phi18*/	4,0,2,2,1,1,3,98,0,2,98,2,7,
/* out0376_em-eta16-phi18*/	3,0,1,1,0,2,4,98,0,6,
/* out0377_em-eta17-phi18*/	4,0,0,4,0,2,2,98,0,3,128,1,2,
/* out0378_em-eta18-phi18*/	2,0,0,3,128,1,4,
/* out0379_em-eta19-phi18*/	2,128,0,2,128,1,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	1,144,3,2,
/* out0382_em-eta2-phi19*/	2,144,2,11,144,3,14,
/* out0383_em-eta3-phi19*/	2,143,3,13,144,2,5,
/* out0384_em-eta4-phi19*/	6,22,1,9,22,2,6,24,0,1,24,1,2,143,2,13,143,3,3,
/* out0385_em-eta5-phi19*/	8,21,0,6,21,1,3,21,2,14,22,0,8,22,1,7,24,1,5,142,3,15,143,2,3,
/* out0386_em-eta6-phi19*/	8,17,1,3,17,2,3,20,0,2,20,2,4,21,0,7,21,1,7,142,2,15,142,3,1,
/* out0387_em-eta7-phi19*/	6,16,2,6,17,1,5,20,0,11,141,4,1,141,5,16,142,2,1,
/* out0388_em-eta8-phi19*/	5,16,0,2,16,1,10,16,2,6,141,3,1,141,4,15,
/* out0389_em-eta9-phi19*/	5,15,0,3,15,2,8,16,0,1,16,1,4,141,3,15,
/* out0390_em-eta10-phi19*/	3,15,0,11,15,1,1,140,3,14,
/* out0391_em-eta11-phi19*/	9,2,1,3,2,2,4,14,0,1,15,0,1,15,1,1,100,0,10,100,2,3,140,2,16,140,3,2,
/* out0392_em-eta12-phi19*/	6,1,2,1,2,1,6,14,0,2,99,2,2,100,1,1,100,2,12,
/* out0393_em-eta13-phi19*/	3,1,2,7,99,0,4,99,2,7,
/* out0394_em-eta14-phi19*/	5,1,0,2,1,1,3,1,2,1,99,0,7,99,1,2,
/* out0395_em-eta15-phi19*/	7,1,0,2,1,1,3,98,0,2,98,2,1,99,1,1,129,1,3,129,2,2,
/* out0396_em-eta16-phi19*/	4,0,2,4,7,1,1,98,0,3,129,1,3,
/* out0397_em-eta17-phi19*/	3,0,2,4,128,1,4,128,2,2,
/* out0398_em-eta18-phi19*/	3,0,0,2,128,0,1,128,1,4,
/* out0399_em-eta19-phi19*/	1,128,0,5,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	1,149,0,2,
/* out0402_em-eta2-phi20*/	2,149,0,14,149,1,11,
/* out0403_em-eta3-phi20*/	2,148,0,13,149,1,5,
/* out0404_em-eta4-phi20*/	4,22,0,1,22,2,10,148,0,3,148,1,13,
/* out0405_em-eta5-phi20*/	7,18,0,2,18,1,10,18,2,14,21,0,2,22,0,7,147,0,15,148,1,3,
/* out0406_em-eta6-phi20*/	8,17,0,5,17,1,1,17,2,13,18,0,1,18,1,6,21,0,1,147,0,1,147,1,15,
/* out0407_em-eta7-phi20*/	8,4,1,1,4,2,3,16,2,3,17,0,8,17,1,7,146,0,16,146,1,1,147,1,1,
/* out0408_em-eta8-phi20*/	6,3,2,1,4,1,5,16,0,11,16,2,1,146,1,15,146,2,1,
/* out0409_em-eta9-phi20*/	4,3,1,5,3,2,8,16,0,2,146,2,15,
/* out0410_em-eta10-phi20*/	4,2,2,3,3,1,8,15,0,1,145,0,14,
/* out0411_em-eta11-phi20*/	8,2,0,2,2,1,1,2,2,8,100,0,6,100,1,6,131,1,2,145,0,2,145,1,16,
/* out0412_em-eta12-phi20*/	5,2,0,4,2,1,5,100,1,9,100,2,1,130,2,3,
/* out0413_em-eta13-phi20*/	7,1,0,2,1,2,3,2,1,1,8,1,1,99,0,3,130,1,6,130,2,2,
/* out0414_em-eta14-phi20*/	4,1,0,6,99,0,2,129,2,5,130,1,3,
/* out0415_em-eta15-phi20*/	4,1,0,3,7,2,2,129,1,2,129,2,5,
/* out0416_em-eta16-phi20*/	3,7,1,2,7,2,2,129,1,6,
/* out0417_em-eta17-phi20*/	3,7,1,4,128,2,5,129,1,1,
/* out0418_em-eta18-phi20*/	3,7,1,1,128,0,2,128,2,4,
/* out0419_em-eta19-phi20*/	1,128,0,4,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	1,149,3,2,
/* out0422_em-eta2-phi21*/	2,149,2,11,149,3,14,
/* out0423_em-eta3-phi21*/	2,148,3,13,149,2,5,
/* out0424_em-eta4-phi21*/	3,6,2,5,148,2,13,148,3,3,
/* out0425_em-eta5-phi21*/	7,5,2,2,6,1,12,6,2,4,18,0,11,18,2,2,147,3,15,148,2,3,
/* out0426_em-eta6-phi21*/	7,5,0,2,5,1,10,5,2,11,17,0,1,18,0,2,147,2,15,147,3,1,
/* out0427_em-eta7-phi21*/	7,4,0,2,4,2,13,5,1,5,17,0,2,146,4,1,146,5,16,147,2,1,
/* out0428_em-eta8-phi21*/	5,3,2,1,4,0,6,4,1,10,146,3,1,146,4,15,
/* out0429_em-eta9-phi21*/	4,3,0,8,3,2,6,10,1,1,146,3,15,
/* out0430_em-eta10-phi21*/	4,3,0,7,3,1,3,9,2,3,145,3,14,
/* out0431_em-eta11-phi21*/	7,2,0,5,2,2,1,9,1,4,131,0,5,131,1,7,145,2,16,145,3,2,
/* out0432_em-eta12-phi21*/	4,2,0,5,8,2,3,130,2,8,131,1,7,
/* out0433_em-eta13-phi21*/	5,8,1,4,8,2,4,130,0,5,130,1,3,130,2,3,
/* out0434_em-eta14-phi21*/	5,1,0,1,8,1,5,129,2,3,130,0,2,130,1,4,
/* out0435_em-eta15-phi21*/	3,7,2,5,129,0,7,129,2,1,
/* out0436_em-eta16-phi21*/	3,7,1,1,7,2,3,129,0,6,
/* out0437_em-eta17-phi21*/	6,7,1,4,95,1,2,95,2,2,128,2,1,129,0,1,129,1,1,
/* out0438_em-eta18-phi21*/	3,7,1,2,95,1,2,128,2,3,
/* out0439_em-eta19-phi21*/	2,128,0,2,128,2,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	1,154,0,2,
/* out0442_em-eta2-phi22*/	2,154,0,14,154,1,11,
/* out0443_em-eta3-phi22*/	2,153,0,13,154,1,5,
/* out0444_em-eta4-phi22*/	6,6,0,2,6,2,5,13,0,1,13,1,3,153,0,3,153,1,13,
/* out0445_em-eta5-phi22*/	8,5,2,1,6,0,14,6,1,4,6,2,2,12,2,8,13,1,4,152,0,15,153,1,3,
/* out0446_em-eta6-phi22*/	6,5,0,12,5,2,2,11,2,3,12,1,9,152,0,1,152,1,15,
/* out0447_em-eta7-phi22*/	8,4,0,3,5,0,2,5,1,1,11,1,9,11,2,7,151,0,16,151,1,1,152,1,1,
/* out0448_em-eta8-phi22*/	5,4,0,5,10,2,11,11,1,3,151,1,15,151,2,1,
/* out0449_em-eta9-phi22*/	4,3,0,1,10,1,12,10,2,2,151,2,15,
/* out0450_em-eta10-phi22*/	3,9,2,11,10,1,1,150,0,14,
/* out0451_em-eta11-phi22*/	7,9,0,2,9,1,8,9,2,1,97,2,1,131,0,7,150,0,2,150,1,16,
/* out0452_em-eta12-phi22*/	6,8,2,6,9,1,3,97,1,4,97,2,5,130,0,2,131,0,4,
/* out0453_em-eta13-phi22*/	6,8,0,3,8,1,1,8,2,3,96,2,2,97,1,4,130,0,6,
/* out0454_em-eta14-phi22*/	5,8,0,2,8,1,4,96,1,2,96,2,7,130,0,1,
/* out0455_em-eta15-phi22*/	5,7,0,1,7,2,3,8,1,1,96,1,7,129,0,1,
/* out0456_em-eta16-phi22*/	5,7,0,4,7,2,1,95,2,5,96,1,1,129,0,1,
/* out0457_em-eta17-phi22*/	3,7,0,3,95,1,2,95,2,4,
/* out0458_em-eta18-phi22*/	3,7,0,1,7,1,1,95,1,5,
/* out0459_em-eta19-phi22*/	1,95,1,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	1,154,3,2,
/* out0462_em-eta2-phi23*/	2,154,2,11,154,3,14,
/* out0463_em-eta3-phi23*/	2,153,3,13,154,2,5,
/* out0464_em-eta4-phi23*/	4,13,0,9,13,1,1,153,2,13,153,3,3,
/* out0465_em-eta5-phi23*/	6,12,0,7,12,2,8,13,0,6,13,1,8,152,3,15,153,2,3,
/* out0466_em-eta6-phi23*/	6,11,0,1,11,2,3,12,0,9,12,1,7,152,2,15,152,3,1,
/* out0467_em-eta7-phi23*/	6,11,0,14,11,1,2,11,2,3,151,4,1,151,5,16,152,2,1,
/* out0468_em-eta8-phi23*/	6,10,0,5,10,2,3,11,0,1,11,1,2,151,3,1,151,4,15,
/* out0469_em-eta9-phi23*/	3,10,0,11,10,1,1,151,3,15,
/* out0470_em-eta10-phi23*/	4,9,0,5,9,2,1,10,1,1,150,3,14,
/* out0471_em-eta11-phi23*/	5,9,0,8,97,0,1,97,2,5,150,2,16,150,3,2,
/* out0472_em-eta12-phi23*/	6,8,0,2,9,0,1,9,1,1,97,0,13,97,1,2,97,2,5,
/* out0473_em-eta13-phi23*/	5,8,0,6,96,0,1,96,2,3,97,0,2,97,1,6,
/* out0474_em-eta14-phi23*/	3,8,0,3,96,0,5,96,2,4,
/* out0475_em-eta15-phi23*/	3,7,0,1,96,0,4,96,1,5,
/* out0476_em-eta16-phi23*/	5,7,0,3,95,0,7,95,2,4,96,0,6,96,1,1,
/* out0477_em-eta17-phi23*/	3,7,0,3,95,0,5,95,2,1,
/* out0478_em-eta18-phi23*/	2,95,0,3,95,1,2,
/* out0479_em-eta19-phi23*/	2,95,0,1,95,1,2
};