parameter integer matrixH [0:2186] = {
/* num inputs = 155(in0-in154) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 5 */
//* total number of input in adders 853 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	1, 99, 6, 
/* out0003_had-eta3-phi0*/	2, 98, 3, 99, 2, 
/* out0004_had-eta4-phi0*/	3, 87, 1, 94, 2, 98, 4, 
/* out0005_had-eta5-phi0*/	3, 94, 12, 97, 4, 98, 1, 
/* out0006_had-eta6-phi0*/	3, 93, 10, 94, 1, 97, 4, 
/* out0007_had-eta7-phi0*/	3, 92, 4, 93, 5, 96, 3, 
/* out0008_had-eta8-phi0*/	2, 92, 7, 96, 3, 
/* out0009_had-eta9-phi0*/	3, 91, 5, 92, 1, 96, 2, 
/* out0010_had-eta10-phi0*/	2, 91, 5, 95, 6, 
/* out0011_had-eta11-phi0*/	3, 90, 3, 91, 1, 95, 2, 
/* out0012_had-eta12-phi0*/	1, 90, 4, 
/* out0013_had-eta13-phi0*/	2, 89, 1, 90, 2, 
/* out0014_had-eta14-phi0*/	1, 89, 2, 
/* out0015_had-eta15-phi0*/	1, 89, 2, 
/* out0016_had-eta16-phi0*/	1, 89, 2, 
/* out0017_had-eta17-phi0*/	1, 88, 3, 
/* out0018_had-eta18-phi0*/	1, 88, 2, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	1, 99, 6, 
/* out0023_had-eta3-phi1*/	2, 98, 3, 99, 2, 
/* out0024_had-eta4-phi1*/	2, 87, 7, 98, 4, 
/* out0025_had-eta5-phi1*/	5, 86, 7, 87, 7, 94, 1, 97, 4, 98, 1, 
/* out0026_had-eta6-phi1*/	4, 85, 2, 86, 5, 93, 1, 97, 4, 
/* out0027_had-eta7-phi1*/	3, 85, 7, 92, 1, 96, 3, 
/* out0028_had-eta8-phi1*/	4, 84, 3, 85, 1, 92, 3, 96, 3, 
/* out0029_had-eta9-phi1*/	3, 84, 3, 91, 2, 96, 2, 
/* out0030_had-eta10-phi1*/	3, 83, 2, 91, 3, 95, 6, 
/* out0031_had-eta11-phi1*/	3, 83, 2, 90, 2, 95, 2, 
/* out0032_had-eta12-phi1*/	1, 90, 3, 
/* out0033_had-eta13-phi1*/	3, 82, 1, 89, 1, 90, 2, 
/* out0034_had-eta14-phi1*/	1, 89, 2, 
/* out0035_had-eta15-phi1*/	1, 89, 2, 
/* out0036_had-eta16-phi1*/	2, 88, 1, 89, 2, 
/* out0037_had-eta17-phi1*/	1, 88, 3, 
/* out0038_had-eta18-phi1*/	1, 88, 2, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	1, 104, 6, 
/* out0043_had-eta3-phi2*/	2, 103, 3, 104, 2, 
/* out0044_had-eta4-phi2*/	3, 80, 4, 87, 1, 103, 4, 
/* out0045_had-eta5-phi2*/	5, 79, 1, 80, 9, 86, 2, 102, 4, 103, 1, 
/* out0046_had-eta6-phi2*/	4, 79, 6, 85, 1, 86, 2, 102, 4, 
/* out0047_had-eta7-phi2*/	4, 78, 2, 79, 1, 85, 5, 101, 3, 
/* out0048_had-eta8-phi2*/	3, 78, 1, 84, 5, 101, 3, 
/* out0049_had-eta9-phi2*/	2, 84, 5, 101, 2, 
/* out0050_had-eta10-phi2*/	2, 83, 4, 100, 6, 
/* out0051_had-eta11-phi2*/	2, 83, 4, 100, 2, 
/* out0052_had-eta12-phi2*/	1, 82, 2, 
/* out0053_had-eta13-phi2*/	1, 82, 2, 
/* out0054_had-eta14-phi2*/	2, 82, 1, 89, 1, 
/* out0055_had-eta15-phi2*/	2, 81, 1, 89, 1, 
/* out0056_had-eta16-phi2*/	1, 81, 1, 
/* out0057_had-eta17-phi2*/	1, 88, 2, 
/* out0058_had-eta18-phi2*/	1, 88, 2, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	0, 
/* out0062_had-eta2-phi3*/	1, 104, 6, 
/* out0063_had-eta3-phi3*/	2, 103, 3, 104, 2, 
/* out0064_had-eta4-phi3*/	2, 74, 1, 103, 4, 
/* out0065_had-eta5-phi3*/	5, 74, 7, 79, 2, 80, 3, 102, 4, 103, 1, 
/* out0066_had-eta6-phi3*/	4, 73, 2, 74, 1, 79, 6, 102, 4, 
/* out0067_had-eta7-phi3*/	2, 78, 7, 101, 3, 
/* out0068_had-eta8-phi3*/	3, 77, 1, 78, 4, 101, 3, 
/* out0069_had-eta9-phi3*/	2, 77, 5, 101, 2, 
/* out0070_had-eta10-phi3*/	3, 77, 1, 83, 2, 100, 6, 
/* out0071_had-eta11-phi3*/	3, 76, 1, 83, 2, 100, 2, 
/* out0072_had-eta12-phi3*/	1, 82, 3, 
/* out0073_had-eta13-phi3*/	1, 82, 2, 
/* out0074_had-eta14-phi3*/	2, 81, 1, 82, 2, 
/* out0075_had-eta15-phi3*/	1, 81, 2, 
/* out0076_had-eta16-phi3*/	1, 81, 1, 
/* out0077_had-eta17-phi3*/	1, 81, 1, 
/* out0078_had-eta18-phi3*/	1, 88, 1, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	0, 
/* out0082_had-eta2-phi4*/	1, 109, 6, 
/* out0083_had-eta3-phi4*/	2, 108, 3, 109, 2, 
/* out0084_had-eta4-phi4*/	2, 74, 1, 108, 4, 
/* out0085_had-eta5-phi4*/	4, 74, 6, 75, 4, 107, 4, 108, 1, 
/* out0086_had-eta6-phi4*/	2, 73, 9, 107, 4, 
/* out0087_had-eta7-phi4*/	4, 72, 3, 73, 3, 78, 1, 106, 3, 
/* out0088_had-eta8-phi4*/	4, 72, 4, 77, 2, 78, 1, 106, 3, 
/* out0089_had-eta9-phi4*/	2, 77, 5, 106, 2, 
/* out0090_had-eta10-phi4*/	3, 76, 3, 77, 2, 105, 6, 
/* out0091_had-eta11-phi4*/	2, 76, 4, 105, 2, 
/* out0092_had-eta12-phi4*/	2, 76, 2, 82, 1, 
/* out0093_had-eta13-phi4*/	2, 60, 1, 82, 1, 
/* out0094_had-eta14-phi4*/	3, 60, 1, 81, 1, 82, 1, 
/* out0095_had-eta15-phi4*/	1, 81, 2, 
/* out0096_had-eta16-phi4*/	1, 81, 1, 
/* out0097_had-eta17-phi4*/	1, 81, 1, 
/* out0098_had-eta18-phi4*/	0, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	0, 
/* out0102_had-eta2-phi5*/	1, 109, 6, 
/* out0103_had-eta3-phi5*/	2, 108, 3, 109, 2, 
/* out0104_had-eta4-phi5*/	1, 108, 4, 
/* out0105_had-eta5-phi5*/	3, 75, 10, 107, 4, 108, 1, 
/* out0106_had-eta6-phi5*/	4, 68, 5, 73, 2, 75, 2, 107, 4, 
/* out0107_had-eta7-phi5*/	3, 68, 2, 72, 4, 106, 3, 
/* out0108_had-eta8-phi5*/	3, 66, 1, 72, 5, 106, 3, 
/* out0109_had-eta9-phi5*/	2, 66, 5, 106, 2, 
/* out0110_had-eta10-phi5*/	3, 66, 2, 76, 2, 105, 6, 
/* out0111_had-eta11-phi5*/	2, 76, 3, 105, 2, 
/* out0112_had-eta12-phi5*/	2, 60, 2, 76, 1, 
/* out0113_had-eta13-phi5*/	1, 60, 2, 
/* out0114_had-eta14-phi5*/	1, 60, 2, 
/* out0115_had-eta15-phi5*/	1, 81, 2, 
/* out0116_had-eta16-phi5*/	1, 81, 1, 
/* out0117_had-eta17-phi5*/	1, 81, 1, 
/* out0118_had-eta18-phi5*/	0, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	0, 
/* out0122_had-eta2-phi6*/	1, 114, 6, 
/* out0123_had-eta3-phi6*/	2, 113, 3, 114, 2, 
/* out0124_had-eta4-phi6*/	1, 113, 4, 
/* out0125_had-eta5-phi6*/	3, 70, 10, 112, 4, 113, 1, 
/* out0126_had-eta6-phi6*/	4, 68, 6, 69, 2, 70, 2, 112, 4, 
/* out0127_had-eta7-phi6*/	3, 67, 4, 68, 3, 111, 3, 
/* out0128_had-eta8-phi6*/	3, 66, 1, 67, 5, 111, 3, 
/* out0129_had-eta9-phi6*/	2, 66, 5, 111, 2, 
/* out0130_had-eta10-phi6*/	3, 61, 2, 66, 2, 110, 6, 
/* out0131_had-eta11-phi6*/	2, 61, 3, 110, 2, 
/* out0132_had-eta12-phi6*/	2, 60, 2, 61, 1, 
/* out0133_had-eta13-phi6*/	1, 60, 2, 
/* out0134_had-eta14-phi6*/	1, 60, 2, 
/* out0135_had-eta15-phi6*/	1, 53, 2, 
/* out0136_had-eta16-phi6*/	1, 53, 1, 
/* out0137_had-eta17-phi6*/	1, 53, 1, 
/* out0138_had-eta18-phi6*/	0, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	0, 
/* out0142_had-eta2-phi7*/	1, 114, 6, 
/* out0143_had-eta3-phi7*/	2, 113, 3, 114, 2, 
/* out0144_had-eta4-phi7*/	2, 71, 1, 113, 4, 
/* out0145_had-eta5-phi7*/	4, 70, 4, 71, 6, 112, 4, 113, 1, 
/* out0146_had-eta6-phi7*/	2, 69, 9, 112, 4, 
/* out0147_had-eta7-phi7*/	4, 63, 1, 67, 3, 69, 3, 111, 3, 
/* out0148_had-eta8-phi7*/	4, 62, 2, 63, 1, 67, 4, 111, 3, 
/* out0149_had-eta9-phi7*/	2, 62, 5, 111, 2, 
/* out0150_had-eta10-phi7*/	3, 61, 3, 62, 1, 110, 6, 
/* out0151_had-eta11-phi7*/	2, 61, 4, 110, 2, 
/* out0152_had-eta12-phi7*/	2, 54, 1, 61, 2, 
/* out0153_had-eta13-phi7*/	2, 54, 1, 60, 1, 
/* out0154_had-eta14-phi7*/	3, 53, 1, 54, 1, 60, 1, 
/* out0155_had-eta15-phi7*/	1, 53, 2, 
/* out0156_had-eta16-phi7*/	1, 53, 1, 
/* out0157_had-eta17-phi7*/	1, 53, 1, 
/* out0158_had-eta18-phi7*/	0, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	0, 
/* out0162_had-eta2-phi8*/	1, 119, 6, 
/* out0163_had-eta3-phi8*/	2, 118, 3, 119, 2, 
/* out0164_had-eta4-phi8*/	2, 71, 1, 118, 4, 
/* out0165_had-eta5-phi8*/	5, 64, 2, 65, 3, 71, 7, 117, 4, 118, 1, 
/* out0166_had-eta6-phi8*/	4, 64, 6, 69, 2, 71, 1, 117, 4, 
/* out0167_had-eta7-phi8*/	2, 63, 7, 116, 3, 
/* out0168_had-eta8-phi8*/	3, 62, 2, 63, 4, 116, 3, 
/* out0169_had-eta9-phi8*/	2, 62, 5, 116, 2, 
/* out0170_had-eta10-phi8*/	3, 55, 2, 62, 1, 115, 6, 
/* out0171_had-eta11-phi8*/	3, 55, 2, 61, 1, 115, 2, 
/* out0172_had-eta12-phi8*/	1, 54, 3, 
/* out0173_had-eta13-phi8*/	1, 54, 2, 
/* out0174_had-eta14-phi8*/	2, 53, 1, 54, 2, 
/* out0175_had-eta15-phi8*/	1, 53, 2, 
/* out0176_had-eta16-phi8*/	1, 53, 1, 
/* out0177_had-eta17-phi8*/	1, 53, 1, 
/* out0178_had-eta18-phi8*/	1, 46, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	0, 
/* out0182_had-eta2-phi9*/	1, 119, 6, 
/* out0183_had-eta3-phi9*/	2, 118, 3, 119, 2, 
/* out0184_had-eta4-phi9*/	3, 59, 1, 65, 4, 118, 4, 
/* out0185_had-eta5-phi9*/	5, 58, 2, 64, 1, 65, 9, 117, 4, 118, 1, 
/* out0186_had-eta6-phi9*/	4, 57, 1, 58, 2, 64, 6, 117, 4, 
/* out0187_had-eta7-phi9*/	4, 57, 5, 63, 2, 64, 1, 116, 3, 
/* out0188_had-eta8-phi9*/	3, 56, 5, 63, 1, 116, 3, 
/* out0189_had-eta9-phi9*/	2, 56, 5, 116, 2, 
/* out0190_had-eta10-phi9*/	2, 55, 4, 115, 6, 
/* out0191_had-eta11-phi9*/	2, 55, 4, 115, 2, 
/* out0192_had-eta12-phi9*/	1, 54, 2, 
/* out0193_had-eta13-phi9*/	1, 54, 2, 
/* out0194_had-eta14-phi9*/	2, 47, 1, 54, 1, 
/* out0195_had-eta15-phi9*/	2, 47, 1, 53, 1, 
/* out0196_had-eta16-phi9*/	1, 53, 1, 
/* out0197_had-eta17-phi9*/	1, 46, 2, 
/* out0198_had-eta18-phi9*/	1, 46, 2, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	0, 
/* out0202_had-eta2-phi10*/	1, 124, 6, 
/* out0203_had-eta3-phi10*/	2, 123, 3, 124, 2, 
/* out0204_had-eta4-phi10*/	2, 59, 7, 123, 4, 
/* out0205_had-eta5-phi10*/	5, 52, 1, 58, 7, 59, 7, 122, 4, 123, 1, 
/* out0206_had-eta6-phi10*/	4, 51, 1, 57, 2, 58, 5, 122, 4, 
/* out0207_had-eta7-phi10*/	3, 50, 1, 57, 7, 121, 3, 
/* out0208_had-eta8-phi10*/	4, 50, 2, 56, 3, 57, 1, 121, 3, 
/* out0209_had-eta9-phi10*/	3, 49, 2, 56, 3, 121, 2, 
/* out0210_had-eta10-phi10*/	3, 49, 2, 55, 2, 120, 6, 
/* out0211_had-eta11-phi10*/	3, 48, 2, 55, 2, 120, 2, 
/* out0212_had-eta12-phi10*/	1, 48, 3, 
/* out0213_had-eta13-phi10*/	3, 47, 1, 48, 1, 54, 1, 
/* out0214_had-eta14-phi10*/	1, 47, 2, 
/* out0215_had-eta15-phi10*/	1, 47, 2, 
/* out0216_had-eta16-phi10*/	1, 47, 1, 
/* out0217_had-eta17-phi10*/	1, 46, 2, 
/* out0218_had-eta18-phi10*/	1, 46, 2, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	0, 
/* out0222_had-eta2-phi11*/	1, 124, 6, 
/* out0223_had-eta3-phi11*/	2, 123, 3, 124, 2, 
/* out0224_had-eta4-phi11*/	3, 52, 2, 59, 1, 123, 4, 
/* out0225_had-eta5-phi11*/	3, 52, 10, 122, 4, 123, 1, 
/* out0226_had-eta6-phi11*/	3, 51, 8, 52, 1, 122, 4, 
/* out0227_had-eta7-phi11*/	3, 50, 3, 51, 4, 121, 3, 
/* out0228_had-eta8-phi11*/	2, 50, 6, 121, 3, 
/* out0229_had-eta9-phi11*/	3, 49, 4, 50, 1, 121, 2, 
/* out0230_had-eta10-phi11*/	2, 49, 4, 120, 6, 
/* out0231_had-eta11-phi11*/	3, 48, 3, 49, 1, 120, 2, 
/* out0232_had-eta12-phi11*/	1, 48, 3, 
/* out0233_had-eta13-phi11*/	2, 47, 1, 48, 2, 
/* out0234_had-eta14-phi11*/	1, 47, 2, 
/* out0235_had-eta15-phi11*/	1, 47, 2, 
/* out0236_had-eta16-phi11*/	1, 47, 1, 
/* out0237_had-eta17-phi11*/	1, 46, 2, 
/* out0238_had-eta18-phi11*/	1, 46, 2, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	0, 
/* out0242_had-eta2-phi12*/	1, 129, 6, 
/* out0243_had-eta3-phi12*/	2, 128, 3, 129, 2, 
/* out0244_had-eta4-phi12*/	2, 45, 5, 128, 4, 
/* out0245_had-eta5-phi12*/	5, 44, 5, 45, 7, 52, 2, 127, 4, 128, 1, 
/* out0246_had-eta6-phi12*/	4, 43, 1, 44, 5, 51, 2, 127, 4, 
/* out0247_had-eta7-phi12*/	4, 43, 6, 50, 1, 51, 1, 126, 3, 
/* out0248_had-eta8-phi12*/	4, 42, 3, 43, 1, 50, 2, 126, 3, 
/* out0249_had-eta9-phi12*/	3, 42, 4, 49, 1, 126, 2, 
/* out0250_had-eta10-phi12*/	3, 41, 2, 49, 2, 125, 6, 
/* out0251_had-eta11-phi12*/	2, 41, 3, 125, 2, 
/* out0252_had-eta12-phi12*/	2, 40, 1, 48, 2, 
/* out0253_had-eta13-phi12*/	1, 40, 2, 
/* out0254_had-eta14-phi12*/	2, 40, 1, 47, 1, 
/* out0255_had-eta15-phi12*/	1, 47, 1, 
/* out0256_had-eta16-phi12*/	1, 39, 1, 
/* out0257_had-eta17-phi12*/	2, 39, 1, 46, 1, 
/* out0258_had-eta18-phi12*/	1, 46, 2, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	0, 
/* out0262_had-eta2-phi13*/	1, 129, 6, 
/* out0263_had-eta3-phi13*/	2, 128, 3, 129, 2, 
/* out0264_had-eta4-phi13*/	3, 38, 2, 45, 2, 128, 4, 
/* out0265_had-eta5-phi13*/	5, 38, 7, 44, 3, 45, 2, 127, 4, 128, 1, 
/* out0266_had-eta6-phi13*/	4, 37, 4, 43, 1, 44, 3, 127, 4, 
/* out0267_had-eta7-phi13*/	4, 36, 1, 37, 1, 43, 6, 126, 3, 
/* out0268_had-eta8-phi13*/	4, 36, 1, 42, 4, 43, 1, 126, 3, 
/* out0269_had-eta9-phi13*/	2, 42, 5, 126, 2, 
/* out0270_had-eta10-phi13*/	2, 41, 4, 125, 6, 
/* out0271_had-eta11-phi13*/	2, 41, 4, 125, 2, 
/* out0272_had-eta12-phi13*/	2, 40, 2, 41, 1, 
/* out0273_had-eta13-phi13*/	1, 40, 3, 
/* out0274_had-eta14-phi13*/	1, 40, 2, 
/* out0275_had-eta15-phi13*/	1, 39, 2, 
/* out0276_had-eta16-phi13*/	1, 39, 1, 
/* out0277_had-eta17-phi13*/	1, 39, 1, 
/* out0278_had-eta18-phi13*/	1, 39, 1, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	0, 
/* out0282_had-eta2-phi14*/	1, 134, 6, 
/* out0283_had-eta3-phi14*/	2, 133, 3, 134, 2, 
/* out0284_had-eta4-phi14*/	2, 38, 2, 133, 4, 
/* out0285_had-eta5-phi14*/	5, 32, 4, 37, 1, 38, 5, 132, 4, 133, 1, 
/* out0286_had-eta6-phi14*/	3, 32, 1, 37, 8, 132, 4, 
/* out0287_had-eta7-phi14*/	4, 31, 1, 36, 5, 37, 2, 131, 3, 
/* out0288_had-eta8-phi14*/	2, 36, 6, 131, 3, 
/* out0289_had-eta9-phi14*/	2, 35, 5, 131, 2, 
/* out0290_had-eta10-phi14*/	3, 35, 3, 41, 1, 130, 6, 
/* out0291_had-eta11-phi14*/	3, 34, 2, 41, 1, 130, 2, 
/* out0292_had-eta12-phi14*/	2, 34, 2, 40, 1, 
/* out0293_had-eta13-phi14*/	1, 40, 2, 
/* out0294_had-eta14-phi14*/	1, 40, 2, 
/* out0295_had-eta15-phi14*/	1, 39, 2, 
/* out0296_had-eta16-phi14*/	1, 39, 1, 
/* out0297_had-eta17-phi14*/	1, 39, 1, 
/* out0298_had-eta18-phi14*/	1, 39, 1, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	0, 
/* out0302_had-eta2-phi15*/	1, 134, 6, 
/* out0303_had-eta3-phi15*/	2, 133, 3, 134, 2, 
/* out0304_had-eta4-phi15*/	2, 28, 5, 133, 4, 
/* out0305_had-eta5-phi15*/	5, 26, 1, 28, 3, 32, 9, 132, 4, 133, 1, 
/* out0306_had-eta6-phi15*/	3, 31, 6, 32, 2, 132, 4, 
/* out0307_had-eta7-phi15*/	4, 30, 1, 31, 5, 36, 1, 131, 3, 
/* out0308_had-eta8-phi15*/	4, 30, 4, 35, 1, 36, 2, 131, 3, 
/* out0309_had-eta9-phi15*/	3, 30, 1, 35, 4, 131, 2, 
/* out0310_had-eta10-phi15*/	3, 34, 1, 35, 3, 130, 6, 
/* out0311_had-eta11-phi15*/	2, 34, 4, 130, 2, 
/* out0312_had-eta12-phi15*/	1, 34, 3, 
/* out0313_had-eta13-phi15*/	1, 33, 2, 
/* out0314_had-eta14-phi15*/	1, 33, 2, 
/* out0315_had-eta15-phi15*/	2, 33, 1, 39, 1, 
/* out0316_had-eta16-phi15*/	1, 39, 1, 
/* out0317_had-eta17-phi15*/	1, 39, 1, 
/* out0318_had-eta18-phi15*/	1, 39, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	0, 
/* out0322_had-eta2-phi16*/	1, 139, 6, 
/* out0323_had-eta3-phi16*/	2, 138, 3, 139, 2, 
/* out0324_had-eta4-phi16*/	3, 27, 1, 28, 4, 138, 4, 
/* out0325_had-eta5-phi16*/	5, 26, 8, 27, 2, 28, 4, 137, 4, 138, 1, 
/* out0326_had-eta6-phi16*/	4, 25, 2, 26, 5, 31, 2, 137, 4, 
/* out0327_had-eta7-phi16*/	4, 25, 4, 30, 2, 31, 2, 136, 3, 
/* out0328_had-eta8-phi16*/	2, 30, 6, 136, 3, 
/* out0329_had-eta9-phi16*/	3, 29, 4, 30, 2, 136, 2, 
/* out0330_had-eta10-phi16*/	2, 29, 4, 135, 6, 
/* out0331_had-eta11-phi16*/	3, 29, 1, 34, 2, 135, 2, 
/* out0332_had-eta12-phi16*/	2, 14, 1, 34, 2, 
/* out0333_had-eta13-phi16*/	1, 33, 2, 
/* out0334_had-eta14-phi16*/	1, 33, 2, 
/* out0335_had-eta15-phi16*/	1, 33, 2, 
/* out0336_had-eta16-phi16*/	1, 0, 1, 
/* out0337_had-eta17-phi16*/	1, 0, 1, 
/* out0338_had-eta18-phi16*/	1, 0, 1, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	0, 
/* out0342_had-eta2-phi17*/	1, 139, 6, 
/* out0343_had-eta3-phi17*/	2, 138, 3, 139, 2, 
/* out0344_had-eta4-phi17*/	2, 27, 4, 138, 4, 
/* out0345_had-eta5-phi17*/	5, 23, 4, 26, 1, 27, 9, 137, 4, 138, 1, 
/* out0346_had-eta6-phi17*/	4, 23, 4, 25, 4, 26, 1, 137, 4, 
/* out0347_had-eta7-phi17*/	3, 19, 1, 25, 6, 136, 3, 
/* out0348_had-eta8-phi17*/	2, 19, 5, 136, 3, 
/* out0349_had-eta9-phi17*/	3, 19, 2, 29, 3, 136, 2, 
/* out0350_had-eta10-phi17*/	2, 29, 4, 135, 6, 
/* out0351_had-eta11-phi17*/	2, 14, 3, 135, 2, 
/* out0352_had-eta12-phi17*/	1, 14, 3, 
/* out0353_had-eta13-phi17*/	2, 14, 1, 33, 2, 
/* out0354_had-eta14-phi17*/	1, 33, 2, 
/* out0355_had-eta15-phi17*/	2, 0, 1, 33, 1, 
/* out0356_had-eta16-phi17*/	1, 0, 2, 
/* out0357_had-eta17-phi17*/	1, 0, 1, 
/* out0358_had-eta18-phi17*/	1, 0, 1, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	0, 
/* out0362_had-eta2-phi18*/	1, 144, 6, 
/* out0363_had-eta3-phi18*/	2, 143, 3, 144, 2, 
/* out0364_had-eta4-phi18*/	2, 24, 4, 143, 4, 
/* out0365_had-eta5-phi18*/	5, 21, 1, 23, 4, 24, 9, 142, 4, 143, 1, 
/* out0366_had-eta6-phi18*/	4, 20, 4, 21, 1, 23, 4, 142, 4, 
/* out0367_had-eta7-phi18*/	3, 19, 1, 20, 6, 141, 3, 
/* out0368_had-eta8-phi18*/	2, 19, 5, 141, 3, 
/* out0369_had-eta9-phi18*/	3, 15, 3, 19, 2, 141, 2, 
/* out0370_had-eta10-phi18*/	2, 15, 4, 140, 6, 
/* out0371_had-eta11-phi18*/	2, 14, 3, 140, 2, 
/* out0372_had-eta12-phi18*/	1, 14, 3, 
/* out0373_had-eta13-phi18*/	2, 1, 2, 14, 1, 
/* out0374_had-eta14-phi18*/	1, 1, 2, 
/* out0375_had-eta15-phi18*/	2, 0, 1, 1, 1, 
/* out0376_had-eta16-phi18*/	1, 0, 2, 
/* out0377_had-eta17-phi18*/	1, 0, 1, 
/* out0378_had-eta18-phi18*/	1, 0, 1, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	0, 
/* out0382_had-eta2-phi19*/	1, 144, 6, 
/* out0383_had-eta3-phi19*/	2, 143, 3, 144, 2, 
/* out0384_had-eta4-phi19*/	3, 22, 4, 24, 1, 143, 4, 
/* out0385_had-eta5-phi19*/	5, 21, 8, 22, 4, 24, 2, 142, 4, 143, 1, 
/* out0386_had-eta6-phi19*/	4, 17, 2, 20, 2, 21, 5, 142, 4, 
/* out0387_had-eta7-phi19*/	4, 16, 2, 17, 2, 20, 4, 141, 3, 
/* out0388_had-eta8-phi19*/	2, 16, 6, 141, 3, 
/* out0389_had-eta9-phi19*/	3, 15, 4, 16, 2, 141, 2, 
/* out0390_had-eta10-phi19*/	2, 15, 4, 140, 6, 
/* out0391_had-eta11-phi19*/	3, 2, 2, 15, 1, 140, 2, 
/* out0392_had-eta12-phi19*/	2, 2, 2, 14, 1, 
/* out0393_had-eta13-phi19*/	1, 1, 2, 
/* out0394_had-eta14-phi19*/	1, 1, 2, 
/* out0395_had-eta15-phi19*/	1, 1, 2, 
/* out0396_had-eta16-phi19*/	1, 0, 1, 
/* out0397_had-eta17-phi19*/	1, 0, 1, 
/* out0398_had-eta18-phi19*/	1, 0, 1, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	0, 
/* out0402_had-eta2-phi20*/	1, 149, 6, 
/* out0403_had-eta3-phi20*/	2, 148, 3, 149, 2, 
/* out0404_had-eta4-phi20*/	2, 22, 5, 148, 4, 
/* out0405_had-eta5-phi20*/	5, 18, 9, 21, 1, 22, 3, 147, 4, 148, 1, 
/* out0406_had-eta6-phi20*/	3, 17, 6, 18, 2, 147, 4, 
/* out0407_had-eta7-phi20*/	4, 4, 1, 16, 1, 17, 5, 146, 3, 
/* out0408_had-eta8-phi20*/	4, 3, 1, 4, 2, 16, 4, 146, 3, 
/* out0409_had-eta9-phi20*/	3, 3, 4, 16, 1, 146, 2, 
/* out0410_had-eta10-phi20*/	3, 2, 1, 3, 3, 145, 6, 
/* out0411_had-eta11-phi20*/	2, 2, 4, 145, 2, 
/* out0412_had-eta12-phi20*/	1, 2, 3, 
/* out0413_had-eta13-phi20*/	1, 1, 2, 
/* out0414_had-eta14-phi20*/	1, 1, 2, 
/* out0415_had-eta15-phi20*/	2, 1, 1, 7, 1, 
/* out0416_had-eta16-phi20*/	1, 7, 1, 
/* out0417_had-eta17-phi20*/	1, 7, 1, 
/* out0418_had-eta18-phi20*/	1, 7, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	0, 
/* out0422_had-eta2-phi21*/	1, 149, 6, 
/* out0423_had-eta3-phi21*/	2, 148, 3, 149, 2, 
/* out0424_had-eta4-phi21*/	2, 6, 2, 148, 4, 
/* out0425_had-eta5-phi21*/	5, 5, 1, 6, 5, 18, 4, 147, 4, 148, 1, 
/* out0426_had-eta6-phi21*/	3, 5, 8, 18, 1, 147, 4, 
/* out0427_had-eta7-phi21*/	4, 4, 5, 5, 2, 17, 1, 146, 3, 
/* out0428_had-eta8-phi21*/	2, 4, 6, 146, 3, 
/* out0429_had-eta9-phi21*/	2, 3, 5, 146, 2, 
/* out0430_had-eta10-phi21*/	3, 3, 3, 9, 1, 145, 6, 
/* out0431_had-eta11-phi21*/	3, 2, 2, 9, 1, 145, 2, 
/* out0432_had-eta12-phi21*/	2, 2, 2, 8, 1, 
/* out0433_had-eta13-phi21*/	1, 8, 2, 
/* out0434_had-eta14-phi21*/	1, 8, 2, 
/* out0435_had-eta15-phi21*/	1, 7, 2, 
/* out0436_had-eta16-phi21*/	1, 7, 1, 
/* out0437_had-eta17-phi21*/	1, 7, 1, 
/* out0438_had-eta18-phi21*/	1, 7, 1, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	0, 
/* out0442_had-eta2-phi22*/	1, 154, 6, 
/* out0443_had-eta3-phi22*/	2, 153, 3, 154, 2, 
/* out0444_had-eta4-phi22*/	3, 6, 2, 13, 2, 153, 4, 
/* out0445_had-eta5-phi22*/	5, 6, 7, 12, 3, 13, 2, 152, 4, 153, 1, 
/* out0446_had-eta6-phi22*/	4, 5, 4, 11, 1, 12, 3, 152, 4, 
/* out0447_had-eta7-phi22*/	4, 4, 1, 5, 1, 11, 6, 151, 3, 
/* out0448_had-eta8-phi22*/	4, 4, 1, 10, 4, 11, 1, 151, 3, 
/* out0449_had-eta9-phi22*/	2, 10, 5, 151, 2, 
/* out0450_had-eta10-phi22*/	2, 9, 4, 150, 6, 
/* out0451_had-eta11-phi22*/	2, 9, 4, 150, 2, 
/* out0452_had-eta12-phi22*/	2, 8, 2, 9, 1, 
/* out0453_had-eta13-phi22*/	1, 8, 3, 
/* out0454_had-eta14-phi22*/	1, 8, 2, 
/* out0455_had-eta15-phi22*/	1, 7, 2, 
/* out0456_had-eta16-phi22*/	1, 7, 1, 
/* out0457_had-eta17-phi22*/	1, 7, 1, 
/* out0458_had-eta18-phi22*/	1, 7, 1, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	0, 
/* out0462_had-eta2-phi23*/	1, 154, 6, 
/* out0463_had-eta3-phi23*/	2, 153, 3, 154, 2, 
/* out0464_had-eta4-phi23*/	2, 13, 5, 153, 4, 
/* out0465_had-eta5-phi23*/	4, 12, 5, 13, 7, 152, 4, 153, 1, 
/* out0466_had-eta6-phi23*/	3, 11, 1, 12, 5, 152, 4, 
/* out0467_had-eta7-phi23*/	2, 11, 6, 151, 3, 
/* out0468_had-eta8-phi23*/	3, 10, 3, 11, 1, 151, 3, 
/* out0469_had-eta9-phi23*/	2, 10, 4, 151, 2, 
/* out0470_had-eta10-phi23*/	2, 9, 2, 150, 6, 
/* out0471_had-eta11-phi23*/	2, 9, 3, 150, 2, 
/* out0472_had-eta12-phi23*/	1, 8, 1, 
/* out0473_had-eta13-phi23*/	1, 8, 2, 
/* out0474_had-eta14-phi23*/	1, 8, 1, 
/* out0475_had-eta15-phi23*/	0, 
/* out0476_had-eta16-phi23*/	1, 7, 1, 
/* out0477_had-eta17-phi23*/	1, 7, 1, 
/* out0478_had-eta18-phi23*/	0, 
/* out0479_had-eta19-phi23*/	0, 
};