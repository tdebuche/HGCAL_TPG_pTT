parameter integer matrixH [0:6087] = {
/* num inputs = 160(in0-in159) */
/* num outputs = 480(out0-out479 */
//* max inputs per outputs = 10 */
//* total number of input in adders 1869 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	1, 137, 0, 3, 
/* out0002_had-eta2-phi0*/	2, 39, 1, 6, 137, 0, 4, 
/* out0003_had-eta3-phi0*/	6, 28, 2, 13, 38, 1, 3, 38, 2, 11, 39, 1, 7, 136, 0, 4, 137, 0, 1, 
/* out0004_had-eta4-phi0*/	6, 28, 0, 16, 28, 1, 4, 28, 2, 3, 37, 2, 8, 38, 1, 7, 136, 0, 4, 
/* out0005_had-eta5-phi0*/	7, 27, 0, 13, 27, 1, 1, 27, 2, 16, 28, 1, 12, 36, 2, 2, 37, 1, 8, 37, 2, 1, 
/* out0006_had-eta6-phi0*/	6, 26, 0, 5, 26, 2, 4, 27, 0, 3, 27, 1, 15, 36, 1, 5, 36, 2, 5, 
/* out0007_had-eta7-phi0*/	5, 25, 2, 11, 26, 0, 11, 26, 1, 5, 26, 2, 12, 35, 2, 4, 
/* out0008_had-eta8-phi0*/	5, 25, 0, 10, 25, 1, 11, 25, 2, 5, 26, 1, 11, 35, 1, 3, 
/* out0009_had-eta9-phi0*/	5, 24, 2, 2, 25, 0, 6, 25, 1, 5, 34, 1, 1, 34, 2, 2, 
/* out0010_had-eta10-phi0*/	3, 24, 0, 8, 24, 1, 11, 24, 2, 14, 
/* out0011_had-eta11-phi0*/	3, 9, 11, 2, 24, 0, 6, 24, 1, 4, 
/* out0012_had-eta12-phi0*/	7, 3, 2, 2, 3, 3, 12, 3, 8, 16, 3, 9, 16, 3, 10, 3, 9, 5, 2, 24, 1, 1, 
/* out0013_had-eta13-phi0*/	6, 3, 0, 1, 3, 1, 5, 3, 2, 14, 3, 3, 2, 3, 6, 4, 3, 10, 13, 
/* out0014_had-eta14-phi0*/	6, 1, 8, 16, 1, 9, 6, 3, 1, 6, 3, 4, 16, 3, 6, 12, 3, 7, 16, 
/* out0015_had-eta15-phi0*/	4, 1, 2, 1, 1, 3, 6, 1, 9, 10, 1, 10, 3, 
/* out0016_had-eta16-phi0*/	4, 1, 2, 12, 1, 3, 1, 1, 6, 1, 1, 10, 13, 
/* out0017_had-eta17-phi0*/	4, 1, 1, 3, 1, 2, 3, 1, 6, 15, 1, 7, 7, 
/* out0018_had-eta18-phi0*/	4, 0, 3, 16, 0, 4, 4, 1, 4, 16, 1, 7, 8, 
/* out0019_had-eta19-phi0*/	4, 0, 1, 16, 0, 2, 1, 0, 4, 8, 0, 5, 16, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	1, 137, 0, 3, 
/* out0022_had-eta2-phi1*/	3, 39, 0, 11, 51, 2, 7, 137, 0, 4, 
/* out0023_had-eta3-phi1*/	10, 38, 0, 12, 38, 1, 1, 38, 2, 5, 39, 0, 5, 39, 1, 3, 50, 2, 3, 51, 1, 12, 51, 2, 7, 136, 0, 4, 137, 0, 1, 
/* out0024_had-eta4-phi1*/	7, 37, 0, 8, 37, 2, 7, 38, 0, 4, 38, 1, 5, 50, 1, 7, 50, 2, 6, 136, 0, 4, 
/* out0025_had-eta5-phi1*/	6, 36, 0, 2, 36, 2, 5, 37, 0, 8, 37, 1, 8, 49, 1, 2, 49, 2, 4, 
/* out0026_had-eta6-phi1*/	3, 36, 0, 12, 36, 1, 9, 36, 2, 4, 
/* out0027_had-eta7-phi1*/	4, 35, 0, 6, 35, 1, 1, 35, 2, 12, 36, 1, 2, 
/* out0028_had-eta8-phi1*/	3, 34, 2, 3, 35, 0, 2, 35, 1, 12, 
/* out0029_had-eta9-phi1*/	3, 34, 0, 1, 34, 1, 3, 34, 2, 10, 
/* out0030_had-eta10-phi1*/	4, 9, 8, 6, 9, 9, 1, 24, 0, 1, 34, 1, 9, 
/* out0031_had-eta11-phi1*/	6, 9, 6, 1, 9, 8, 10, 9, 9, 2, 9, 10, 9, 9, 11, 14, 24, 0, 1, 
/* out0032_had-eta12-phi1*/	5, 3, 0, 2, 3, 3, 2, 9, 4, 9, 9, 5, 14, 9, 6, 6, 
/* out0033_had-eta13-phi1*/	4, 3, 0, 13, 3, 1, 2, 8, 8, 10, 9, 4, 3, 
/* out0034_had-eta14-phi1*/	3, 3, 1, 3, 8, 5, 5, 8, 11, 15, 
/* out0035_had-eta15-phi1*/	4, 1, 0, 2, 1, 3, 7, 8, 4, 3, 8, 5, 8, 
/* out0036_had-eta16-phi1*/	3, 1, 0, 11, 1, 1, 2, 1, 3, 2, 
/* out0037_had-eta17-phi1*/	4, 1, 0, 2, 1, 1, 9, 2, 8, 1, 2, 11, 2, 
/* out0038_had-eta18-phi1*/	6, 0, 2, 4, 0, 4, 3, 1, 1, 2, 1, 7, 1, 2, 5, 3, 2, 11, 4, 
/* out0039_had-eta19-phi1*/	3, 0, 2, 10, 0, 4, 1, 2, 5, 1, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	1, 139, 0, 3, 
/* out0042_had-eta2-phi2*/	5, 51, 0, 4, 51, 2, 2, 63, 0, 3, 63, 1, 14, 139, 0, 4, 
/* out0043_had-eta3-phi2*/	9, 50, 0, 3, 50, 2, 4, 51, 0, 12, 51, 1, 4, 62, 1, 8, 62, 2, 13, 63, 1, 1, 138, 0, 4, 139, 0, 1, 
/* out0044_had-eta4-phi2*/	9, 49, 0, 1, 49, 2, 3, 50, 0, 13, 50, 1, 9, 50, 2, 3, 61, 1, 2, 61, 2, 5, 62, 1, 1, 138, 0, 4, 
/* out0045_had-eta5-phi2*/	3, 49, 0, 12, 49, 1, 10, 49, 2, 9, 
/* out0046_had-eta6-phi2*/	5, 36, 0, 2, 48, 0, 3, 48, 1, 1, 48, 2, 16, 49, 1, 4, 
/* out0047_had-eta7-phi2*/	3, 35, 0, 5, 47, 2, 4, 48, 1, 12, 
/* out0048_had-eta8-phi2*/	5, 34, 0, 1, 34, 2, 1, 35, 0, 3, 47, 1, 5, 47, 2, 7, 
/* out0049_had-eta9-phi2*/	3, 34, 0, 11, 46, 2, 1, 47, 1, 2, 
/* out0050_had-eta10-phi2*/	6, 9, 3, 4, 9, 9, 8, 34, 0, 3, 34, 1, 3, 46, 1, 1, 46, 2, 2, 
/* out0051_had-eta11-phi2*/	7, 9, 0, 1, 9, 1, 1, 9, 2, 13, 9, 3, 12, 9, 6, 1, 9, 9, 5, 9, 10, 7, 
/* out0052_had-eta12-phi2*/	5, 9, 1, 6, 9, 2, 3, 9, 4, 2, 9, 6, 8, 9, 7, 14, 
/* out0053_had-eta13-phi2*/	5, 8, 8, 6, 8, 9, 14, 8, 10, 4, 9, 4, 2, 9, 7, 1, 
/* out0054_had-eta14-phi2*/	4, 8, 2, 2, 8, 6, 8, 8, 10, 12, 8, 11, 1, 
/* out0055_had-eta15-phi2*/	4, 8, 4, 7, 8, 5, 3, 8, 6, 6, 8, 7, 3, 
/* out0056_had-eta16-phi2*/	3, 1, 0, 1, 2, 8, 10, 8, 4, 5, 
/* out0057_had-eta17-phi2*/	3, 2, 8, 4, 2, 10, 2, 2, 11, 7, 
/* out0058_had-eta18-phi2*/	4, 2, 5, 6, 2, 6, 1, 2, 10, 1, 2, 11, 3, 
/* out0059_had-eta19-phi2*/	4, 0, 0, 16, 0, 2, 1, 2, 4, 3, 2, 5, 5, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 139, 0, 3, 
/* out0062_had-eta2-phi3*/	6, 63, 0, 13, 63, 1, 1, 123, 0, 4, 123, 1, 6, 123, 2, 16, 139, 0, 4, 
/* out0063_had-eta3-phi3*/	8, 62, 0, 16, 62, 1, 6, 62, 2, 3, 121, 1, 2, 121, 2, 9, 123, 1, 8, 138, 0, 4, 139, 0, 1, 
/* out0064_had-eta4-phi3*/	6, 61, 0, 15, 61, 1, 8, 61, 2, 11, 62, 1, 1, 121, 1, 2, 138, 0, 4, 
/* out0065_had-eta5-phi3*/	5, 49, 0, 3, 60, 0, 3, 60, 1, 2, 60, 2, 16, 61, 1, 6, 
/* out0066_had-eta6-phi3*/	3, 48, 0, 10, 59, 2, 4, 60, 1, 11, 
/* out0067_had-eta7-phi3*/	6, 47, 0, 4, 47, 2, 3, 48, 0, 3, 48, 1, 3, 59, 1, 4, 59, 2, 4, 
/* out0068_had-eta8-phi3*/	3, 47, 0, 10, 47, 1, 5, 47, 2, 2, 
/* out0069_had-eta9-phi3*/	3, 46, 0, 1, 46, 2, 9, 47, 1, 4, 
/* out0070_had-eta10-phi3*/	3, 46, 0, 1, 46, 1, 7, 46, 2, 4, 
/* out0071_had-eta11-phi3*/	3, 9, 0, 14, 10, 8, 10, 46, 1, 4, 
/* out0072_had-eta12-phi3*/	6, 9, 0, 1, 9, 1, 9, 9, 7, 1, 10, 5, 4, 10, 8, 2, 10, 11, 15, 
/* out0073_had-eta13-phi3*/	6, 8, 0, 3, 8, 2, 1, 8, 3, 14, 8, 9, 2, 10, 4, 1, 10, 5, 6, 
/* out0074_had-eta14-phi3*/	4, 8, 0, 4, 8, 1, 5, 8, 2, 12, 8, 3, 2, 
/* out0075_had-eta15-phi3*/	4, 8, 1, 5, 8, 2, 1, 8, 6, 2, 8, 7, 12, 
/* out0076_had-eta16-phi3*/	4, 2, 8, 1, 2, 9, 13, 8, 4, 1, 8, 7, 1, 
/* out0077_had-eta17-phi3*/	3, 2, 2, 2, 2, 9, 1, 2, 10, 11, 
/* out0078_had-eta18-phi3*/	2, 2, 6, 9, 2, 10, 2, 
/* out0079_had-eta19-phi3*/	4, 2, 4, 12, 2, 5, 1, 2, 6, 2, 2, 7, 1, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 141, 0, 3, 
/* out0082_had-eta2-phi4*/	5, 123, 0, 11, 124, 0, 2, 124, 1, 1, 124, 2, 15, 141, 0, 4, 
/* out0083_had-eta3-phi4*/	10, 121, 0, 15, 121, 1, 4, 121, 2, 7, 122, 2, 4, 123, 0, 1, 123, 1, 2, 124, 1, 11, 124, 2, 1, 140, 0, 4, 141, 0, 1, 
/* out0084_had-eta4-phi4*/	9, 61, 0, 1, 120, 0, 8, 120, 1, 2, 120, 2, 16, 121, 0, 1, 121, 1, 8, 122, 1, 1, 122, 2, 1, 140, 0, 4, 
/* out0085_had-eta5-phi4*/	3, 60, 0, 11, 119, 2, 7, 120, 1, 12, 
/* out0086_had-eta6-phi4*/	6, 59, 0, 7, 59, 2, 6, 60, 0, 2, 60, 1, 3, 119, 1, 4, 119, 2, 3, 
/* out0087_had-eta7-phi4*/	4, 58, 2, 1, 59, 0, 6, 59, 1, 12, 59, 2, 2, 
/* out0088_had-eta8-phi4*/	3, 47, 0, 2, 58, 1, 1, 58, 2, 13, 
/* out0089_had-eta9-phi4*/	2, 46, 0, 6, 58, 1, 7, 
/* out0090_had-eta10-phi4*/	3, 46, 0, 8, 46, 1, 2, 70, 2, 1, 
/* out0091_had-eta11-phi4*/	6, 10, 2, 2, 10, 3, 6, 10, 8, 4, 10, 9, 16, 10, 10, 4, 46, 1, 2, 
/* out0092_had-eta12-phi4*/	5, 10, 2, 6, 10, 5, 1, 10, 6, 13, 10, 10, 12, 10, 11, 1, 
/* out0093_had-eta13-phi4*/	6, 8, 0, 2, 10, 4, 14, 10, 5, 5, 10, 6, 2, 10, 7, 3, 14, 8, 1, 
/* out0094_had-eta14-phi4*/	4, 8, 0, 7, 8, 1, 2, 14, 8, 9, 14, 11, 3, 
/* out0095_had-eta15-phi4*/	4, 2, 9, 1, 8, 1, 4, 14, 5, 4, 14, 11, 9, 
/* out0096_had-eta16-phi4*/	3, 2, 3, 12, 2, 9, 1, 14, 5, 2, 
/* out0097_had-eta17-phi4*/	3, 2, 1, 1, 2, 2, 9, 2, 3, 4, 
/* out0098_had-eta18-phi4*/	4, 2, 1, 2, 2, 2, 5, 2, 6, 4, 2, 7, 1, 
/* out0099_had-eta19-phi4*/	2, 2, 4, 1, 2, 7, 9, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 141, 0, 3, 
/* out0102_had-eta2-phi5*/	2, 124, 0, 11, 141, 0, 4, 
/* out0103_had-eta3-phi5*/	7, 122, 0, 15, 122, 1, 2, 122, 2, 11, 124, 0, 3, 124, 1, 4, 140, 0, 4, 141, 0, 1, 
/* out0104_had-eta4-phi5*/	5, 120, 0, 7, 122, 0, 1, 122, 1, 13, 130, 2, 14, 140, 0, 4, 
/* out0105_had-eta5-phi5*/	6, 119, 0, 12, 119, 2, 6, 120, 0, 1, 120, 1, 2, 130, 1, 7, 130, 2, 2, 
/* out0106_had-eta6-phi5*/	4, 59, 0, 1, 119, 0, 4, 119, 1, 12, 125, 2, 7, 
/* out0107_had-eta7-phi5*/	5, 58, 0, 1, 58, 2, 1, 59, 0, 2, 125, 1, 7, 125, 2, 9, 
/* out0108_had-eta8-phi5*/	4, 58, 0, 14, 58, 1, 1, 58, 2, 1, 125, 1, 1, 
/* out0109_had-eta9-phi5*/	3, 58, 0, 1, 58, 1, 7, 70, 2, 6, 
/* out0110_had-eta10-phi5*/	2, 70, 1, 3, 70, 2, 9, 
/* out0111_had-eta11-phi5*/	3, 10, 0, 9, 10, 3, 9, 70, 1, 5, 
/* out0112_had-eta12-phi5*/	6, 10, 0, 7, 10, 1, 14, 10, 2, 8, 10, 3, 1, 10, 6, 1, 10, 7, 1, 
/* out0113_had-eta13-phi5*/	5, 10, 1, 2, 10, 4, 1, 10, 7, 12, 14, 8, 2, 14, 9, 9, 
/* out0114_had-eta14-phi5*/	4, 14, 8, 4, 14, 9, 6, 14, 10, 11, 14, 11, 2, 
/* out0115_had-eta15-phi5*/	4, 14, 5, 6, 14, 6, 7, 14, 10, 4, 14, 11, 2, 
/* out0116_had-eta16-phi5*/	3, 2, 0, 4, 14, 4, 7, 14, 5, 4, 
/* out0117_had-eta17-phi5*/	2, 2, 0, 11, 2, 1, 1, 
/* out0118_had-eta18-phi5*/	2, 2, 0, 1, 2, 1, 10, 
/* out0119_had-eta19-phi5*/	2, 2, 1, 2, 2, 7, 5, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 143, 0, 3, 
/* out0122_had-eta2-phi6*/	2, 132, 2, 11, 143, 0, 4, 
/* out0123_had-eta3-phi6*/	7, 131, 0, 11, 131, 1, 2, 131, 2, 15, 132, 1, 4, 132, 2, 3, 142, 0, 4, 143, 0, 1, 
/* out0124_had-eta4-phi6*/	6, 127, 2, 7, 130, 0, 14, 130, 1, 1, 131, 1, 13, 131, 2, 1, 142, 0, 4, 
/* out0125_had-eta5-phi6*/	6, 126, 0, 6, 126, 2, 12, 127, 1, 2, 127, 2, 1, 130, 0, 2, 130, 1, 8, 
/* out0126_had-eta6-phi6*/	4, 72, 2, 1, 125, 0, 7, 126, 1, 12, 126, 2, 4, 
/* out0127_had-eta7-phi6*/	5, 71, 0, 1, 71, 2, 1, 72, 2, 2, 125, 0, 9, 125, 1, 7, 
/* out0128_had-eta8-phi6*/	4, 71, 0, 1, 71, 1, 1, 71, 2, 14, 125, 1, 1, 
/* out0129_had-eta9-phi6*/	3, 70, 0, 6, 71, 1, 7, 71, 2, 1, 
/* out0130_had-eta10-phi6*/	2, 70, 0, 9, 70, 1, 3, 
/* out0131_had-eta11-phi6*/	3, 15, 8, 9, 15, 9, 9, 70, 1, 5, 
/* out0132_had-eta12-phi6*/	6, 15, 5, 1, 15, 6, 1, 15, 8, 7, 15, 9, 1, 15, 10, 8, 15, 11, 14, 
/* out0133_had-eta13-phi6*/	6, 14, 0, 2, 14, 3, 10, 14, 9, 1, 15, 4, 1, 15, 5, 12, 15, 11, 2, 
/* out0134_had-eta14-phi6*/	5, 14, 0, 3, 14, 1, 1, 14, 2, 12, 14, 3, 6, 14, 10, 1, 
/* out0135_had-eta15-phi6*/	4, 14, 1, 1, 14, 2, 4, 14, 6, 9, 14, 7, 5, 
/* out0136_had-eta16-phi6*/	3, 14, 4, 9, 14, 7, 4, 18, 8, 4, 
/* out0137_had-eta17-phi6*/	2, 18, 8, 11, 18, 11, 1, 
/* out0138_had-eta18-phi6*/	2, 18, 8, 1, 18, 11, 10, 
/* out0139_had-eta19-phi6*/	2, 18, 5, 5, 18, 11, 2, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 143, 0, 3, 
/* out0142_had-eta2-phi7*/	5, 129, 2, 11, 132, 0, 15, 132, 1, 1, 132, 2, 2, 143, 0, 4, 
/* out0143_had-eta3-phi7*/	10, 128, 0, 7, 128, 1, 4, 128, 2, 15, 129, 1, 2, 129, 2, 1, 131, 0, 4, 132, 0, 1, 132, 1, 11, 142, 0, 4, 143, 0, 1, 
/* out0144_had-eta4-phi7*/	9, 74, 2, 1, 127, 0, 16, 127, 1, 2, 127, 2, 8, 128, 1, 8, 128, 2, 1, 131, 0, 1, 131, 1, 1, 142, 0, 4, 
/* out0145_had-eta5-phi7*/	3, 73, 2, 11, 126, 0, 7, 127, 1, 12, 
/* out0146_had-eta6-phi7*/	6, 72, 0, 6, 72, 2, 7, 73, 1, 3, 73, 2, 2, 126, 0, 3, 126, 1, 4, 
/* out0147_had-eta7-phi7*/	4, 71, 0, 1, 72, 0, 2, 72, 1, 12, 72, 2, 6, 
/* out0148_had-eta8-phi7*/	3, 71, 0, 13, 71, 1, 1, 85, 2, 2, 
/* out0149_had-eta9-phi7*/	2, 71, 1, 7, 84, 2, 6, 
/* out0150_had-eta10-phi7*/	3, 70, 0, 1, 84, 1, 2, 84, 2, 8, 
/* out0151_had-eta11-phi7*/	6, 15, 0, 4, 15, 2, 4, 15, 3, 16, 15, 9, 6, 15, 10, 2, 84, 1, 2, 
/* out0152_had-eta12-phi7*/	5, 15, 1, 1, 15, 2, 12, 15, 6, 13, 15, 7, 1, 15, 10, 6, 
/* out0153_had-eta13-phi7*/	6, 14, 0, 1, 15, 4, 14, 15, 5, 3, 15, 6, 2, 15, 7, 4, 19, 8, 2, 
/* out0154_had-eta14-phi7*/	4, 14, 0, 10, 14, 1, 4, 19, 8, 7, 19, 11, 2, 
/* out0155_had-eta15-phi7*/	5, 14, 1, 10, 14, 7, 5, 18, 3, 1, 18, 9, 1, 19, 11, 4, 
/* out0156_had-eta16-phi7*/	3, 14, 7, 2, 18, 3, 1, 18, 9, 12, 
/* out0157_had-eta17-phi7*/	3, 18, 9, 3, 18, 10, 9, 18, 11, 1, 
/* out0158_had-eta18-phi7*/	4, 18, 5, 1, 18, 6, 4, 18, 10, 5, 18, 11, 2, 
/* out0159_had-eta19-phi7*/	2, 18, 4, 1, 18, 5, 9, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 145, 0, 3, 
/* out0162_had-eta2-phi8*/	6, 76, 0, 1, 76, 1, 13, 129, 0, 16, 129, 1, 6, 129, 2, 4, 145, 0, 4, 
/* out0163_had-eta3-phi8*/	8, 75, 0, 3, 75, 1, 6, 75, 2, 16, 128, 0, 9, 128, 1, 2, 129, 1, 8, 144, 0, 4, 145, 0, 1, 
/* out0164_had-eta4-phi8*/	6, 74, 0, 11, 74, 1, 8, 74, 2, 15, 75, 1, 1, 128, 1, 2, 144, 0, 4, 
/* out0165_had-eta5-phi8*/	5, 73, 0, 16, 73, 1, 2, 73, 2, 3, 74, 1, 6, 87, 2, 3, 
/* out0166_had-eta6-phi8*/	3, 72, 0, 4, 73, 1, 11, 86, 2, 10, 
/* out0167_had-eta7-phi8*/	6, 72, 0, 4, 72, 1, 4, 85, 0, 3, 85, 2, 4, 86, 1, 3, 86, 2, 3, 
/* out0168_had-eta8-phi8*/	3, 85, 0, 2, 85, 1, 5, 85, 2, 10, 
/* out0169_had-eta9-phi8*/	3, 84, 0, 9, 84, 2, 1, 85, 1, 4, 
/* out0170_had-eta10-phi8*/	3, 84, 0, 4, 84, 1, 7, 84, 2, 1, 
/* out0171_had-eta11-phi8*/	3, 15, 0, 10, 20, 8, 14, 84, 1, 4, 
/* out0172_had-eta12-phi8*/	6, 15, 0, 2, 15, 1, 15, 15, 7, 5, 20, 5, 1, 20, 8, 1, 20, 11, 9, 
/* out0173_had-eta13-phi8*/	6, 15, 4, 1, 15, 7, 6, 19, 3, 2, 19, 8, 3, 19, 9, 15, 19, 10, 1, 
/* out0174_had-eta14-phi8*/	4, 19, 8, 4, 19, 9, 1, 19, 10, 12, 19, 11, 5, 
/* out0175_had-eta15-phi8*/	4, 19, 5, 12, 19, 6, 2, 19, 10, 1, 19, 11, 5, 
/* out0176_had-eta16-phi8*/	4, 18, 0, 1, 18, 3, 13, 19, 4, 1, 19, 5, 1, 
/* out0177_had-eta17-phi8*/	3, 18, 2, 11, 18, 3, 1, 18, 10, 2, 
/* out0178_had-eta18-phi8*/	2, 18, 2, 2, 18, 6, 9, 
/* out0179_had-eta19-phi8*/	4, 18, 4, 12, 18, 5, 1, 18, 6, 2, 18, 7, 1, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 145, 0, 3, 
/* out0182_had-eta2-phi9*/	5, 76, 0, 14, 76, 1, 3, 89, 0, 2, 89, 2, 4, 145, 0, 4, 
/* out0183_had-eta3-phi9*/	9, 75, 0, 13, 75, 1, 8, 76, 0, 1, 88, 0, 4, 88, 2, 3, 89, 1, 4, 89, 2, 12, 144, 0, 4, 145, 0, 1, 
/* out0184_had-eta4-phi9*/	9, 74, 0, 5, 74, 1, 2, 75, 1, 1, 87, 0, 3, 87, 2, 1, 88, 0, 3, 88, 1, 9, 88, 2, 13, 144, 0, 4, 
/* out0185_had-eta5-phi9*/	3, 87, 0, 9, 87, 1, 10, 87, 2, 12, 
/* out0186_had-eta6-phi9*/	5, 86, 0, 16, 86, 1, 1, 86, 2, 3, 87, 1, 4, 98, 2, 2, 
/* out0187_had-eta7-phi9*/	3, 85, 0, 4, 86, 1, 12, 97, 2, 5, 
/* out0188_had-eta8-phi9*/	5, 85, 0, 7, 85, 1, 5, 96, 0, 1, 96, 2, 1, 97, 2, 3, 
/* out0189_had-eta9-phi9*/	3, 84, 0, 1, 85, 1, 2, 96, 2, 11, 
/* out0190_had-eta10-phi9*/	6, 20, 3, 8, 20, 9, 4, 84, 0, 2, 84, 1, 1, 96, 1, 3, 96, 2, 3, 
/* out0191_had-eta11-phi9*/	7, 20, 2, 7, 20, 3, 5, 20, 6, 1, 20, 8, 1, 20, 9, 12, 20, 10, 13, 20, 11, 1, 
/* out0192_had-eta12-phi9*/	5, 20, 4, 2, 20, 5, 14, 20, 6, 8, 20, 10, 3, 20, 11, 6, 
/* out0193_had-eta13-phi9*/	5, 19, 0, 6, 19, 2, 4, 19, 3, 14, 20, 4, 2, 20, 5, 1, 
/* out0194_had-eta14-phi9*/	4, 19, 1, 1, 19, 2, 12, 19, 6, 8, 19, 10, 2, 
/* out0195_had-eta15-phi9*/	4, 19, 4, 7, 19, 5, 3, 19, 6, 6, 19, 7, 3, 
/* out0196_had-eta16-phi9*/	2, 18, 0, 10, 19, 4, 5, 
/* out0197_had-eta17-phi9*/	3, 18, 0, 4, 18, 1, 7, 18, 2, 2, 
/* out0198_had-eta18-phi9*/	4, 18, 1, 3, 18, 2, 1, 18, 6, 1, 18, 7, 6, 
/* out0199_had-eta19-phi9*/	4, 4, 4, 5, 4, 5, 1, 18, 4, 3, 18, 7, 5, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 147, 0, 3, 
/* out0202_had-eta2-phi10*/	3, 89, 0, 7, 101, 1, 11, 147, 0, 4, 
/* out0203_had-eta3-phi10*/	10, 88, 0, 3, 89, 0, 7, 89, 1, 12, 100, 0, 5, 100, 1, 1, 100, 2, 12, 101, 0, 3, 101, 1, 5, 146, 0, 4, 147, 0, 1, 
/* out0204_had-eta4-phi10*/	7, 88, 0, 6, 88, 1, 7, 99, 0, 7, 99, 2, 8, 100, 1, 5, 100, 2, 4, 146, 0, 4, 
/* out0205_had-eta5-phi10*/	6, 87, 0, 4, 87, 1, 2, 98, 0, 5, 98, 2, 2, 99, 1, 8, 99, 2, 8, 
/* out0206_had-eta6-phi10*/	3, 98, 0, 4, 98, 1, 9, 98, 2, 12, 
/* out0207_had-eta7-phi10*/	4, 97, 0, 12, 97, 1, 1, 97, 2, 6, 98, 1, 2, 
/* out0208_had-eta8-phi10*/	3, 96, 0, 3, 97, 1, 12, 97, 2, 2, 
/* out0209_had-eta9-phi10*/	3, 96, 0, 10, 96, 1, 3, 96, 2, 1, 
/* out0210_had-eta10-phi10*/	4, 20, 0, 6, 20, 3, 1, 29, 2, 1, 96, 1, 9, 
/* out0211_had-eta11-phi10*/	6, 20, 0, 10, 20, 1, 14, 20, 2, 9, 20, 3, 2, 20, 6, 1, 29, 2, 1, 
/* out0212_had-eta12-phi10*/	5, 7, 8, 2, 7, 9, 1, 20, 4, 9, 20, 6, 6, 20, 7, 14, 
/* out0213_had-eta13-phi10*/	4, 7, 8, 12, 7, 11, 1, 19, 0, 10, 20, 4, 3, 
/* out0214_had-eta14-phi10*/	3, 7, 11, 3, 19, 1, 15, 19, 7, 5, 
/* out0215_had-eta15-phi10*/	4, 6, 8, 2, 6, 9, 6, 19, 4, 3, 19, 7, 8, 
/* out0216_had-eta16-phi10*/	3, 6, 8, 12, 6, 9, 2, 6, 11, 1, 
/* out0217_had-eta17-phi10*/	4, 6, 8, 2, 6, 11, 8, 18, 0, 1, 18, 1, 2, 
/* out0218_had-eta18-phi10*/	5, 4, 3, 1, 4, 5, 2, 6, 11, 2, 18, 1, 4, 18, 7, 3, 
/* out0219_had-eta19-phi10*/	3, 4, 4, 11, 4, 5, 11, 18, 7, 1, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 147, 0, 3, 
/* out0222_had-eta2-phi11*/	2, 101, 0, 6, 147, 0, 4, 
/* out0223_had-eta3-phi11*/	6, 33, 0, 1, 100, 0, 11, 100, 1, 3, 101, 0, 7, 146, 0, 4, 147, 0, 1, 
/* out0224_had-eta4-phi11*/	6, 33, 0, 2, 33, 1, 3, 33, 2, 16, 99, 0, 8, 100, 1, 7, 146, 0, 4, 
/* out0225_had-eta5-phi11*/	7, 32, 0, 4, 32, 1, 1, 32, 2, 13, 33, 1, 1, 98, 0, 2, 99, 0, 1, 99, 1, 8, 
/* out0226_had-eta6-phi11*/	6, 31, 0, 4, 31, 2, 5, 32, 1, 3, 32, 2, 3, 98, 0, 5, 98, 1, 5, 
/* out0227_had-eta7-phi11*/	3, 31, 1, 4, 31, 2, 11, 97, 0, 4, 
/* out0228_had-eta8-phi11*/	3, 30, 0, 4, 30, 2, 10, 97, 1, 3, 
/* out0229_had-eta9-phi11*/	5, 29, 0, 1, 30, 1, 4, 30, 2, 6, 96, 0, 2, 96, 1, 1, 
/* out0230_had-eta10-phi11*/	2, 29, 0, 3, 29, 2, 8, 
/* out0231_had-eta11-phi11*/	3, 20, 1, 2, 29, 1, 3, 29, 2, 6, 
/* out0232_had-eta12-phi11*/	5, 7, 2, 2, 7, 3, 12, 7, 9, 13, 7, 10, 2, 20, 7, 2, 
/* out0233_had-eta13-phi11*/	6, 7, 2, 1, 7, 6, 3, 7, 8, 2, 7, 9, 2, 7, 10, 14, 7, 11, 5, 
/* out0234_had-eta14-phi11*/	4, 6, 3, 2, 7, 5, 12, 7, 6, 1, 7, 11, 7, 
/* out0235_had-eta15-phi11*/	4, 6, 2, 2, 6, 3, 9, 6, 9, 7, 6, 10, 1, 
/* out0236_had-eta16-phi11*/	5, 6, 2, 2, 6, 6, 1, 6, 9, 1, 6, 10, 12, 6, 11, 1, 
/* out0237_had-eta17-phi11*/	4, 6, 5, 4, 6, 6, 3, 6, 10, 3, 6, 11, 4, 
/* out0238_had-eta18-phi11*/	2, 4, 3, 4, 6, 5, 7, 
/* out0239_had-eta19-phi11*/	4, 4, 2, 2, 4, 3, 7, 4, 5, 2, 4, 6, 16, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 149, 0, 3, 
/* out0242_had-eta2-phi12*/	3, 45, 0, 1, 45, 1, 9, 149, 0, 4, 
/* out0243_had-eta3-phi12*/	7, 33, 0, 2, 44, 0, 4, 44, 2, 11, 45, 0, 4, 45, 1, 7, 148, 0, 4, 149, 0, 1, 
/* out0244_had-eta4-phi12*/	7, 33, 0, 11, 33, 1, 11, 43, 0, 2, 43, 2, 6, 44, 1, 2, 44, 2, 5, 148, 0, 4, 
/* out0245_had-eta5-phi12*/	7, 32, 0, 12, 32, 1, 6, 33, 1, 1, 42, 0, 1, 42, 2, 1, 43, 1, 1, 43, 2, 8, 
/* out0246_had-eta6-phi12*/	3, 31, 0, 9, 32, 1, 6, 42, 2, 10, 
/* out0247_had-eta7-phi12*/	3, 31, 0, 3, 31, 1, 12, 41, 2, 4, 
/* out0248_had-eta8-phi12*/	3, 30, 0, 12, 30, 1, 2, 41, 2, 3, 
/* out0249_had-eta9-phi12*/	3, 29, 0, 1, 30, 1, 10, 40, 2, 3, 
/* out0250_had-eta10-phi12*/	3, 29, 0, 10, 29, 1, 1, 40, 2, 1, 
/* out0251_had-eta11-phi12*/	2, 13, 8, 2, 29, 1, 9, 
/* out0252_had-eta12-phi12*/	6, 7, 0, 15, 7, 1, 5, 7, 2, 5, 7, 3, 4, 13, 8, 2, 29, 1, 1, 
/* out0253_had-eta13-phi12*/	4, 7, 1, 3, 7, 2, 8, 7, 6, 11, 7, 7, 5, 
/* out0254_had-eta14-phi12*/	5, 6, 0, 3, 7, 4, 13, 7, 5, 4, 7, 6, 1, 7, 7, 1, 
/* out0255_had-eta15-phi12*/	4, 6, 0, 9, 6, 1, 2, 6, 2, 3, 6, 3, 5, 
/* out0256_had-eta16-phi12*/	3, 6, 1, 1, 6, 2, 9, 6, 6, 6, 
/* out0257_had-eta17-phi12*/	4, 6, 4, 3, 6, 5, 3, 6, 6, 6, 6, 7, 2, 
/* out0258_had-eta18-phi12*/	3, 4, 0, 3, 6, 4, 6, 6, 5, 2, 
/* out0259_had-eta19-phi12*/	4, 4, 0, 4, 4, 1, 1, 4, 2, 14, 4, 3, 4, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 149, 0, 3, 
/* out0262_had-eta2-phi13*/	4, 45, 0, 6, 57, 0, 5, 57, 2, 2, 149, 0, 4, 
/* out0263_had-eta3-phi13*/	10, 44, 0, 12, 44, 1, 5, 45, 0, 5, 56, 0, 2, 56, 2, 1, 57, 0, 1, 57, 1, 4, 57, 2, 14, 148, 0, 4, 149, 0, 1, 
/* out0264_had-eta4-phi13*/	5, 43, 0, 14, 43, 2, 1, 44, 1, 9, 56, 2, 13, 148, 0, 4, 
/* out0265_had-eta5-phi13*/	4, 42, 0, 8, 43, 1, 15, 43, 2, 1, 55, 2, 6, 
/* out0266_had-eta6-phi13*/	3, 42, 0, 7, 42, 1, 13, 42, 2, 5, 
/* out0267_had-eta7-phi13*/	4, 41, 0, 13, 41, 1, 1, 41, 2, 5, 42, 1, 2, 
/* out0268_had-eta8-phi13*/	3, 40, 0, 3, 41, 1, 9, 41, 2, 4, 
/* out0269_had-eta9-phi13*/	3, 40, 0, 5, 40, 1, 1, 40, 2, 8, 
/* out0270_had-eta10-phi13*/	6, 13, 3, 6, 13, 9, 1, 29, 0, 1, 29, 1, 1, 40, 1, 4, 40, 2, 4, 
/* out0271_had-eta11-phi13*/	6, 13, 2, 2, 13, 3, 6, 13, 8, 6, 13, 9, 15, 13, 10, 8, 29, 1, 1, 
/* out0272_had-eta12-phi13*/	6, 7, 0, 1, 7, 1, 3, 13, 5, 2, 13, 8, 6, 13, 10, 5, 13, 11, 15, 
/* out0273_had-eta13-phi13*/	6, 7, 1, 5, 7, 7, 9, 11, 3, 2, 11, 9, 7, 13, 5, 2, 13, 11, 1, 
/* out0274_had-eta14-phi13*/	6, 7, 4, 3, 7, 7, 1, 11, 8, 12, 11, 9, 7, 11, 10, 1, 11, 11, 1, 
/* out0275_had-eta15-phi13*/	4, 6, 0, 4, 6, 1, 5, 11, 8, 4, 11, 11, 7, 
/* out0276_had-eta16-phi13*/	2, 6, 1, 8, 6, 7, 7, 
/* out0277_had-eta17-phi13*/	4, 5, 8, 2, 5, 9, 1, 6, 4, 4, 6, 7, 6, 
/* out0278_had-eta18-phi13*/	3, 4, 0, 2, 5, 8, 6, 6, 4, 3, 
/* out0279_had-eta19-phi13*/	3, 4, 0, 7, 4, 1, 13, 5, 8, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 151, 0, 3, 
/* out0282_had-eta2-phi14*/	4, 57, 0, 6, 69, 0, 7, 69, 1, 16, 151, 0, 4, 
/* out0283_had-eta3-phi14*/	8, 56, 0, 7, 57, 0, 4, 57, 1, 12, 68, 0, 5, 68, 2, 15, 69, 0, 1, 150, 0, 4, 151, 0, 1, 
/* out0284_had-eta4-phi14*/	9, 55, 0, 4, 56, 0, 7, 56, 1, 16, 56, 2, 2, 67, 0, 1, 67, 2, 7, 68, 1, 1, 68, 2, 1, 150, 0, 4, 
/* out0285_had-eta5-phi14*/	3, 55, 0, 11, 55, 1, 11, 55, 2, 9, 
/* out0286_had-eta6-phi14*/	6, 42, 1, 1, 54, 0, 10, 54, 1, 1, 54, 2, 9, 55, 1, 3, 55, 2, 1, 
/* out0287_had-eta7-phi14*/	6, 41, 0, 3, 41, 1, 2, 53, 0, 2, 53, 2, 1, 54, 1, 5, 54, 2, 7, 
/* out0288_had-eta8-phi14*/	4, 40, 0, 2, 41, 1, 4, 53, 0, 1, 53, 2, 11, 
/* out0289_had-eta9-phi14*/	4, 40, 0, 6, 40, 1, 5, 52, 2, 1, 53, 2, 2, 
/* out0290_had-eta10-phi14*/	4, 13, 0, 11, 13, 3, 1, 40, 1, 6, 52, 2, 3, 
/* out0291_had-eta11-phi14*/	7, 13, 0, 5, 13, 1, 9, 13, 2, 14, 13, 3, 3, 13, 6, 5, 13, 7, 2, 13, 10, 2, 
/* out0292_had-eta12-phi14*/	5, 13, 4, 8, 13, 5, 10, 13, 6, 11, 13, 7, 3, 13, 10, 1, 
/* out0293_had-eta13-phi14*/	6, 11, 0, 6, 11, 2, 4, 11, 3, 14, 11, 9, 1, 13, 4, 1, 13, 5, 2, 
/* out0294_had-eta14-phi14*/	4, 11, 2, 6, 11, 6, 3, 11, 9, 1, 11, 10, 13, 
/* out0295_had-eta15-phi14*/	4, 11, 5, 6, 11, 6, 3, 11, 10, 2, 11, 11, 7, 
/* out0296_had-eta16-phi14*/	5, 5, 3, 6, 5, 9, 3, 6, 7, 1, 11, 5, 4, 11, 11, 1, 
/* out0297_had-eta17-phi14*/	3, 5, 3, 1, 5, 9, 11, 5, 10, 2, 
/* out0298_had-eta18-phi14*/	4, 5, 8, 5, 5, 9, 1, 5, 10, 2, 5, 11, 3, 
/* out0299_had-eta19-phi14*/	3, 4, 1, 2, 5, 8, 2, 5, 11, 7, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 151, 0, 3, 
/* out0302_had-eta2-phi15*/	5, 69, 0, 8, 113, 0, 12, 113, 1, 3, 113, 2, 12, 151, 0, 4, 
/* out0303_had-eta3-phi15*/	8, 68, 0, 11, 68, 1, 14, 111, 0, 2, 111, 2, 9, 113, 1, 4, 113, 2, 4, 150, 0, 4, 151, 0, 1, 
/* out0304_had-eta4-phi15*/	6, 67, 0, 15, 67, 1, 11, 67, 2, 7, 68, 1, 1, 111, 2, 2, 150, 0, 4, 
/* out0305_had-eta5-phi15*/	7, 55, 0, 1, 55, 1, 2, 66, 0, 10, 66, 1, 1, 66, 2, 9, 67, 1, 4, 67, 2, 2, 
/* out0306_had-eta6-phi15*/	6, 54, 0, 6, 54, 1, 4, 65, 0, 2, 65, 2, 2, 66, 1, 4, 66, 2, 7, 
/* out0307_had-eta7-phi15*/	3, 53, 0, 7, 54, 1, 6, 65, 2, 8, 
/* out0308_had-eta8-phi15*/	3, 53, 0, 6, 53, 1, 9, 53, 2, 2, 
/* out0309_had-eta9-phi15*/	3, 52, 0, 8, 52, 2, 2, 53, 1, 5, 
/* out0310_had-eta10-phi15*/	3, 52, 0, 1, 52, 1, 2, 52, 2, 8, 
/* out0311_had-eta11-phi15*/	6, 12, 3, 5, 12, 9, 5, 13, 1, 7, 13, 7, 7, 52, 1, 2, 52, 2, 2, 
/* out0312_had-eta12-phi15*/	5, 12, 8, 12, 12, 9, 10, 12, 11, 1, 13, 4, 7, 13, 7, 4, 
/* out0313_had-eta13-phi15*/	5, 11, 0, 10, 11, 1, 10, 11, 2, 1, 12, 8, 4, 12, 11, 2, 
/* out0314_had-eta14-phi15*/	4, 11, 1, 3, 11, 2, 5, 11, 6, 7, 11, 7, 7, 
/* out0315_had-eta15-phi15*/	4, 11, 4, 11, 11, 5, 5, 11, 6, 3, 11, 7, 1, 
/* out0316_had-eta16-phi15*/	4, 5, 0, 6, 5, 3, 8, 11, 4, 1, 11, 5, 1, 
/* out0317_had-eta17-phi15*/	3, 5, 2, 9, 5, 3, 1, 5, 10, 4, 
/* out0318_had-eta18-phi15*/	3, 5, 6, 3, 5, 10, 8, 5, 11, 1, 
/* out0319_had-eta19-phi15*/	3, 5, 5, 4, 5, 6, 1, 5, 11, 5, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 153, 0, 3, 
/* out0322_had-eta2-phi16*/	6, 112, 0, 11, 112, 1, 1, 112, 2, 7, 113, 0, 4, 113, 1, 6, 153, 0, 4, 
/* out0323_had-eta3-phi16*/	10, 110, 0, 1, 110, 2, 4, 111, 0, 14, 111, 1, 10, 111, 2, 3, 112, 1, 3, 112, 2, 9, 113, 1, 3, 152, 0, 4, 153, 0, 1, 
/* out0324_had-eta4-phi16*/	8, 67, 1, 1, 109, 0, 14, 109, 1, 3, 109, 2, 9, 110, 2, 2, 111, 1, 6, 111, 2, 2, 152, 0, 4, 
/* out0325_had-eta5-phi16*/	6, 66, 0, 6, 66, 1, 5, 108, 0, 3, 108, 2, 4, 109, 1, 5, 109, 2, 7, 
/* out0326_had-eta6-phi16*/	3, 65, 0, 12, 66, 1, 6, 108, 2, 7, 
/* out0327_had-eta7-phi16*/	4, 64, 0, 1, 65, 0, 1, 65, 1, 13, 65, 2, 6, 
/* out0328_had-eta8-phi16*/	3, 53, 1, 2, 64, 0, 6, 64, 2, 9, 
/* out0329_had-eta9-phi16*/	2, 52, 0, 6, 64, 2, 7, 
/* out0330_had-eta10-phi16*/	3, 52, 0, 1, 52, 1, 10, 77, 2, 1, 
/* out0331_had-eta11-phi16*/	5, 12, 0, 13, 12, 1, 1, 12, 2, 5, 12, 3, 11, 52, 1, 2, 
/* out0332_had-eta12-phi16*/	5, 12, 2, 9, 12, 6, 8, 12, 9, 1, 12, 10, 15, 12, 11, 1, 
/* out0333_had-eta13-phi16*/	6, 11, 1, 2, 12, 5, 10, 12, 6, 1, 12, 10, 1, 12, 11, 12, 16, 3, 1, 
/* out0334_had-eta14-phi16*/	4, 11, 1, 1, 11, 7, 8, 16, 3, 2, 16, 9, 10, 
/* out0335_had-eta15-phi16*/	4, 5, 0, 1, 11, 4, 4, 16, 8, 11, 16, 9, 1, 
/* out0336_had-eta16-phi16*/	3, 5, 0, 9, 5, 1, 5, 16, 8, 2, 
/* out0337_had-eta17-phi16*/	4, 5, 1, 4, 5, 2, 7, 5, 6, 3, 5, 7, 1, 
/* out0338_had-eta18-phi16*/	4, 5, 4, 1, 5, 5, 5, 5, 6, 9, 5, 7, 1, 
/* out0339_had-eta19-phi16*/	2, 5, 4, 3, 5, 5, 7, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 153, 0, 3, 
/* out0342_had-eta2-phi17*/	3, 112, 0, 5, 112, 1, 5, 153, 0, 4, 
/* out0343_had-eta3-phi17*/	6, 110, 0, 15, 110, 1, 7, 110, 2, 4, 112, 1, 7, 152, 0, 4, 153, 0, 1, 
/* out0344_had-eta4-phi17*/	7, 109, 0, 2, 109, 1, 5, 110, 1, 9, 110, 2, 6, 133, 0, 8, 133, 2, 7, 152, 0, 4, 
/* out0345_had-eta5-phi17*/	5, 108, 0, 13, 108, 1, 4, 108, 2, 1, 109, 1, 3, 133, 2, 9, 
/* out0346_had-eta6-phi17*/	6, 65, 0, 1, 65, 1, 1, 108, 1, 12, 108, 2, 4, 114, 0, 6, 114, 2, 1, 
/* out0347_had-eta7-phi17*/	4, 64, 0, 1, 65, 1, 2, 114, 0, 2, 114, 2, 14, 
/* out0348_had-eta8-phi17*/	3, 64, 0, 8, 64, 1, 8, 114, 2, 1, 
/* out0349_had-eta9-phi17*/	2, 64, 1, 8, 77, 0, 5, 
/* out0350_had-eta10-phi17*/	2, 77, 0, 2, 77, 2, 10, 
/* out0351_had-eta11-phi17*/	4, 12, 0, 3, 12, 1, 14, 12, 7, 2, 77, 2, 5, 
/* out0352_had-eta12-phi17*/	6, 12, 1, 1, 12, 2, 2, 12, 4, 7, 12, 5, 1, 12, 6, 7, 12, 7, 14, 
/* out0353_had-eta13-phi17*/	4, 12, 4, 9, 12, 5, 5, 16, 0, 7, 16, 3, 4, 
/* out0354_had-eta14-phi17*/	4, 16, 2, 7, 16, 3, 9, 16, 9, 3, 16, 10, 4, 
/* out0355_had-eta15-phi17*/	4, 16, 8, 2, 16, 9, 2, 16, 10, 11, 16, 11, 4, 
/* out0356_had-eta16-phi17*/	3, 5, 1, 3, 16, 8, 1, 16, 11, 11, 
/* out0357_had-eta17-phi17*/	2, 5, 1, 4, 5, 7, 9, 
/* out0358_had-eta18-phi17*/	2, 5, 4, 5, 5, 7, 5, 
/* out0359_had-eta19-phi17*/	1, 5, 4, 7, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 155, 0, 3, 
/* out0362_had-eta2-phi18*/	3, 135, 0, 5, 135, 2, 5, 155, 0, 4, 
/* out0363_had-eta3-phi18*/	6, 134, 0, 15, 134, 1, 4, 134, 2, 7, 135, 2, 7, 154, 0, 4, 155, 0, 1, 
/* out0364_had-eta4-phi18*/	7, 116, 0, 2, 116, 2, 5, 133, 0, 8, 133, 1, 7, 134, 1, 6, 134, 2, 9, 154, 0, 4, 
/* out0365_had-eta5-phi18*/	5, 115, 0, 13, 115, 1, 1, 115, 2, 4, 116, 2, 3, 133, 1, 9, 
/* out0366_had-eta6-phi18*/	6, 79, 0, 1, 79, 2, 1, 114, 0, 6, 114, 1, 1, 115, 1, 4, 115, 2, 12, 
/* out0367_had-eta7-phi18*/	4, 78, 0, 1, 79, 2, 2, 114, 0, 2, 114, 1, 14, 
/* out0368_had-eta8-phi18*/	3, 78, 0, 8, 78, 2, 8, 114, 1, 1, 
/* out0369_had-eta9-phi18*/	2, 77, 0, 6, 78, 2, 8, 
/* out0370_had-eta10-phi18*/	2, 77, 0, 3, 77, 1, 9, 
/* out0371_had-eta11-phi18*/	4, 17, 0, 3, 17, 3, 14, 17, 9, 2, 77, 1, 5, 
/* out0372_had-eta12-phi18*/	6, 17, 2, 2, 17, 3, 1, 17, 8, 7, 17, 9, 14, 17, 10, 7, 17, 11, 1, 
/* out0373_had-eta13-phi18*/	4, 16, 0, 9, 16, 1, 4, 17, 8, 9, 17, 11, 5, 
/* out0374_had-eta14-phi18*/	4, 16, 1, 8, 16, 2, 9, 16, 6, 4, 16, 7, 2, 
/* out0375_had-eta15-phi18*/	5, 16, 4, 1, 16, 5, 5, 16, 6, 12, 16, 7, 1, 16, 10, 1, 
/* out0376_had-eta16-phi18*/	3, 16, 5, 11, 16, 11, 1, 21, 3, 3, 
/* out0377_had-eta17-phi18*/	2, 21, 3, 4, 21, 9, 9, 
/* out0378_had-eta18-phi18*/	2, 21, 8, 5, 21, 9, 5, 
/* out0379_had-eta19-phi18*/	1, 21, 8, 7, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 155, 0, 3, 
/* out0382_had-eta2-phi19*/	6, 118, 0, 4, 118, 2, 6, 135, 0, 11, 135, 1, 7, 135, 2, 1, 155, 0, 4, 
/* out0383_had-eta3-phi19*/	10, 117, 0, 14, 117, 1, 3, 117, 2, 10, 118, 2, 3, 134, 0, 1, 134, 1, 4, 135, 1, 9, 135, 2, 3, 154, 0, 4, 155, 0, 1, 
/* out0384_had-eta4-phi19*/	8, 81, 2, 1, 116, 0, 14, 116, 1, 9, 116, 2, 3, 117, 1, 2, 117, 2, 6, 134, 1, 2, 154, 0, 4, 
/* out0385_had-eta5-phi19*/	6, 80, 0, 6, 80, 2, 5, 115, 0, 3, 115, 1, 4, 116, 1, 7, 116, 2, 5, 
/* out0386_had-eta6-phi19*/	3, 79, 0, 12, 80, 2, 6, 115, 1, 7, 
/* out0387_had-eta7-phi19*/	4, 78, 0, 1, 79, 0, 1, 79, 1, 6, 79, 2, 13, 
/* out0388_had-eta8-phi19*/	3, 78, 0, 6, 78, 1, 9, 91, 2, 2, 
/* out0389_had-eta9-phi19*/	2, 78, 1, 7, 90, 0, 6, 
/* out0390_had-eta10-phi19*/	3, 77, 1, 2, 90, 0, 1, 90, 2, 10, 
/* out0391_had-eta11-phi19*/	5, 17, 0, 13, 17, 1, 11, 17, 2, 5, 17, 3, 1, 90, 2, 2, 
/* out0392_had-eta12-phi19*/	5, 17, 2, 9, 17, 5, 1, 17, 6, 15, 17, 7, 1, 17, 10, 8, 
/* out0393_had-eta13-phi19*/	6, 16, 1, 1, 17, 5, 12, 17, 6, 1, 17, 10, 1, 17, 11, 10, 22, 3, 2, 
/* out0394_had-eta14-phi19*/	4, 16, 1, 3, 16, 7, 11, 22, 3, 1, 22, 9, 8, 
/* out0395_had-eta15-phi19*/	4, 16, 4, 12, 16, 7, 2, 21, 0, 1, 22, 8, 4, 
/* out0396_had-eta16-phi19*/	3, 16, 4, 3, 21, 0, 9, 21, 3, 5, 
/* out0397_had-eta17-phi19*/	4, 21, 2, 7, 21, 3, 4, 21, 9, 1, 21, 10, 3, 
/* out0398_had-eta18-phi19*/	4, 21, 8, 1, 21, 9, 1, 21, 10, 9, 21, 11, 5, 
/* out0399_had-eta19-phi19*/	2, 21, 8, 3, 21, 11, 7, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 157, 0, 3, 
/* out0402_had-eta2-phi20*/	5, 83, 1, 8, 118, 0, 12, 118, 1, 12, 118, 2, 3, 157, 0, 4, 
/* out0403_had-eta3-phi20*/	8, 82, 0, 11, 82, 2, 14, 117, 0, 2, 117, 1, 9, 118, 1, 4, 118, 2, 4, 156, 0, 4, 157, 0, 1, 
/* out0404_had-eta4-phi20*/	6, 81, 0, 15, 81, 1, 7, 81, 2, 11, 82, 2, 1, 117, 1, 2, 156, 0, 4, 
/* out0405_had-eta5-phi20*/	7, 80, 0, 10, 80, 1, 9, 80, 2, 1, 81, 1, 2, 81, 2, 4, 93, 0, 1, 93, 2, 2, 
/* out0406_had-eta6-phi20*/	6, 79, 0, 2, 79, 1, 2, 80, 1, 7, 80, 2, 4, 92, 0, 6, 92, 2, 4, 
/* out0407_had-eta7-phi20*/	3, 79, 1, 8, 91, 0, 7, 92, 2, 6, 
/* out0408_had-eta8-phi20*/	3, 91, 0, 6, 91, 1, 2, 91, 2, 10, 
/* out0409_had-eta9-phi20*/	3, 90, 0, 8, 90, 1, 2, 91, 2, 4, 
/* out0410_had-eta10-phi20*/	3, 90, 0, 1, 90, 1, 8, 90, 2, 2, 
/* out0411_had-eta11-phi20*/	6, 17, 1, 5, 17, 7, 5, 23, 3, 7, 23, 9, 7, 90, 1, 2, 90, 2, 2, 
/* out0412_had-eta12-phi20*/	5, 17, 4, 12, 17, 5, 1, 17, 7, 10, 23, 8, 7, 23, 9, 4, 
/* out0413_had-eta13-phi20*/	5, 17, 4, 4, 17, 5, 2, 22, 0, 10, 22, 2, 1, 22, 3, 10, 
/* out0414_had-eta14-phi20*/	4, 22, 2, 5, 22, 3, 3, 22, 9, 7, 22, 10, 7, 
/* out0415_had-eta15-phi20*/	4, 22, 8, 11, 22, 9, 1, 22, 10, 3, 22, 11, 5, 
/* out0416_had-eta16-phi20*/	4, 21, 0, 6, 21, 1, 8, 22, 8, 1, 22, 11, 1, 
/* out0417_had-eta17-phi20*/	3, 21, 1, 1, 21, 2, 9, 21, 6, 4, 
/* out0418_had-eta18-phi20*/	3, 21, 5, 1, 21, 6, 8, 21, 10, 3, 
/* out0419_had-eta19-phi20*/	3, 21, 5, 5, 21, 10, 1, 21, 11, 4, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 157, 0, 3, 
/* out0422_had-eta2-phi21*/	4, 83, 0, 16, 83, 1, 7, 95, 0, 6, 157, 0, 4, 
/* out0423_had-eta3-phi21*/	8, 82, 0, 5, 82, 1, 15, 83, 1, 1, 94, 0, 7, 95, 0, 4, 95, 2, 12, 156, 0, 4, 157, 0, 1, 
/* out0424_had-eta4-phi21*/	9, 81, 0, 1, 81, 1, 7, 82, 1, 1, 82, 2, 1, 93, 0, 4, 94, 0, 7, 94, 1, 2, 94, 2, 16, 156, 0, 4, 
/* out0425_had-eta5-phi21*/	3, 93, 0, 11, 93, 1, 9, 93, 2, 11, 
/* out0426_had-eta6-phi21*/	6, 92, 0, 10, 92, 1, 9, 92, 2, 1, 93, 1, 1, 93, 2, 3, 104, 2, 1, 
/* out0427_had-eta7-phi21*/	6, 91, 0, 2, 91, 1, 1, 92, 1, 7, 92, 2, 5, 103, 0, 3, 103, 2, 2, 
/* out0428_had-eta8-phi21*/	4, 91, 0, 1, 91, 1, 11, 102, 0, 2, 103, 2, 4, 
/* out0429_had-eta9-phi21*/	4, 90, 1, 1, 91, 1, 2, 102, 0, 6, 102, 2, 5, 
/* out0430_had-eta10-phi21*/	4, 23, 0, 11, 23, 1, 1, 90, 1, 3, 102, 2, 6, 
/* out0431_had-eta11-phi21*/	7, 23, 0, 5, 23, 1, 3, 23, 2, 14, 23, 3, 9, 23, 6, 2, 23, 9, 2, 23, 10, 5, 
/* out0432_had-eta12-phi21*/	5, 23, 6, 1, 23, 8, 8, 23, 9, 3, 23, 10, 11, 23, 11, 10, 
/* out0433_had-eta13-phi21*/	6, 22, 0, 6, 22, 1, 14, 22, 2, 4, 22, 7, 1, 23, 8, 1, 23, 11, 2, 
/* out0434_had-eta14-phi21*/	4, 22, 2, 6, 22, 6, 13, 22, 7, 1, 22, 10, 3, 
/* out0435_had-eta15-phi21*/	4, 22, 5, 7, 22, 6, 2, 22, 10, 3, 22, 11, 6, 
/* out0436_had-eta16-phi21*/	4, 21, 1, 6, 21, 7, 3, 22, 5, 1, 22, 11, 4, 
/* out0437_had-eta17-phi21*/	3, 21, 1, 1, 21, 6, 2, 21, 7, 11, 
/* out0438_had-eta18-phi21*/	4, 21, 4, 5, 21, 5, 3, 21, 6, 2, 21, 7, 1, 
/* out0439_had-eta19-phi21*/	2, 21, 4, 2, 21, 5, 7, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 159, 0, 3, 
/* out0442_had-eta2-phi22*/	4, 95, 0, 5, 95, 1, 2, 107, 1, 6, 159, 0, 4, 
/* out0443_had-eta3-phi22*/	10, 94, 0, 2, 94, 1, 1, 95, 0, 1, 95, 1, 14, 95, 2, 4, 106, 0, 12, 106, 2, 5, 107, 1, 5, 158, 0, 4, 159, 0, 1, 
/* out0444_had-eta4-phi22*/	5, 94, 1, 13, 105, 0, 14, 105, 1, 1, 106, 2, 9, 158, 0, 4, 
/* out0445_had-eta5-phi22*/	4, 93, 1, 6, 104, 0, 8, 105, 1, 1, 105, 2, 15, 
/* out0446_had-eta6-phi22*/	3, 104, 0, 7, 104, 1, 5, 104, 2, 13, 
/* out0447_had-eta7-phi22*/	4, 103, 0, 13, 103, 1, 5, 103, 2, 1, 104, 2, 2, 
/* out0448_had-eta8-phi22*/	3, 102, 0, 3, 103, 1, 4, 103, 2, 9, 
/* out0449_had-eta9-phi22*/	3, 102, 0, 5, 102, 1, 8, 102, 2, 1, 
/* out0450_had-eta10-phi22*/	4, 23, 1, 6, 23, 7, 1, 102, 1, 4, 102, 2, 4, 
/* out0451_had-eta11-phi22*/	5, 23, 1, 6, 23, 2, 2, 23, 4, 6, 23, 6, 8, 23, 7, 15, 
/* out0452_had-eta12-phi22*/	4, 23, 4, 6, 23, 5, 15, 23, 6, 5, 23, 11, 2, 
/* out0453_had-eta13-phi22*/	4, 22, 1, 2, 22, 7, 7, 23, 5, 1, 23, 11, 2, 
/* out0454_had-eta14-phi22*/	4, 22, 4, 12, 22, 5, 1, 22, 6, 1, 22, 7, 7, 
/* out0455_had-eta15-phi22*/	2, 22, 4, 4, 22, 5, 7, 
/* out0456_had-eta16-phi22*/	0, 
/* out0457_had-eta17-phi22*/	2, 21, 4, 2, 21, 7, 1, 
/* out0458_had-eta18-phi22*/	1, 21, 4, 6, 
/* out0459_had-eta19-phi22*/	1, 21, 4, 1, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 159, 0, 3, 
/* out0462_had-eta2-phi23*/	3, 107, 0, 9, 107, 1, 1, 159, 0, 4, 
/* out0463_had-eta3-phi23*/	6, 106, 0, 4, 106, 1, 11, 107, 0, 7, 107, 1, 4, 158, 0, 4, 159, 0, 1, 
/* out0464_had-eta4-phi23*/	5, 105, 0, 2, 105, 1, 6, 106, 1, 5, 106, 2, 2, 158, 0, 4, 
/* out0465_had-eta5-phi23*/	4, 104, 0, 1, 104, 1, 1, 105, 1, 8, 105, 2, 1, 
/* out0466_had-eta6-phi23*/	1, 104, 1, 10, 
/* out0467_had-eta7-phi23*/	1, 103, 1, 4, 
/* out0468_had-eta8-phi23*/	1, 103, 1, 3, 
/* out0469_had-eta9-phi23*/	1, 102, 1, 3, 
/* out0470_had-eta10-phi23*/	1, 102, 1, 1, 
/* out0471_had-eta11-phi23*/	1, 23, 4, 2, 
/* out0472_had-eta12-phi23*/	1, 23, 4, 2, 
/* out0473_had-eta13-phi23*/	0, 
/* out0474_had-eta14-phi23*/	0, 
/* out0475_had-eta15-phi23*/	0, 
/* out0476_had-eta16-phi23*/	0, 
/* out0477_had-eta17-phi23*/	0, 
/* out0478_had-eta18-phi23*/	0, 
/* out0479_had-eta19-phi23*/	0, 
};