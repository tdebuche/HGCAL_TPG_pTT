parameter integer matrixH [0:10536] = {
/* num inputs = 298(in0-in297) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 15 */
//* total number of input in adders 3352 */

/* out0000_had-eta0-phi0*/	1, 253, 0, 1, 
/* out0001_had-eta1-phi0*/	1, 253, 0, 5, 
/* out0002_had-eta2-phi0*/	3, 39, 2, 14, 252, 0, 2, 253, 0, 2, 
/* out0003_had-eta3-phi0*/	3, 38, 2, 10, 39, 1, 12, 252, 0, 4, 
/* out0004_had-eta4-phi0*/	8, 28, 0, 15, 28, 1, 13, 28, 2, 16, 37, 2, 5, 38, 1, 10, 38, 2, 1, 251, 0, 3, 252, 0, 2, 
/* out0005_had-eta5-phi0*/	9, 27, 0, 10, 27, 1, 11, 27, 2, 16, 28, 0, 1, 28, 1, 3, 36, 2, 1, 37, 1, 8, 37, 2, 4, 251, 0, 4, 
/* out0006_had-eta6-phi0*/	8, 26, 0, 3, 26, 2, 4, 27, 0, 6, 27, 1, 5, 36, 1, 4, 36, 2, 6, 250, 0, 2, 251, 0, 1, 
/* out0007_had-eta7-phi0*/	6, 26, 0, 13, 26, 1, 3, 26, 2, 12, 35, 2, 3, 36, 1, 1, 250, 0, 3, 
/* out0008_had-eta8-phi0*/	9, 25, 0, 7, 25, 2, 5, 26, 1, 13, 35, 1, 3, 35, 2, 1, 193, 0, 1, 193, 2, 10, 245, 1, 3, 250, 0, 2, 
/* out0009_had-eta9-phi0*/	11, 24, 2, 10, 25, 0, 9, 25, 1, 5, 25, 2, 11, 34, 2, 2, 193, 0, 6, 193, 1, 7, 193, 2, 6, 244, 2, 4, 245, 1, 9, 250, 0, 1, 
/* out0010_had-eta10-phi0*/	9, 24, 0, 7, 24, 2, 5, 25, 1, 11, 34, 1, 1, 192, 0, 1, 192, 2, 12, 193, 1, 6, 244, 1, 6, 244, 2, 7, 
/* out0011_had-eta11-phi0*/	9, 9, 11, 1, 24, 0, 7, 24, 1, 3, 24, 2, 1, 192, 0, 3, 192, 1, 8, 192, 2, 3, 243, 2, 3, 244, 1, 4, 
/* out0012_had-eta12-phi0*/	11, 3, 3, 10, 3, 8, 16, 3, 9, 16, 3, 10, 2, 9, 5, 2, 9, 11, 2, 24, 1, 13, 191, 2, 7, 192, 1, 5, 243, 1, 4, 243, 2, 5, 
/* out0013_had-eta13-phi0*/	11, 3, 0, 1, 3, 1, 3, 3, 2, 15, 3, 3, 5, 3, 6, 2, 3, 10, 14, 191, 0, 1, 191, 1, 4, 191, 2, 5, 242, 2, 1, 243, 1, 3, 
/* out0014_had-eta14-phi0*/	7, 3, 1, 8, 3, 2, 1, 3, 6, 14, 3, 7, 12, 190, 2, 1, 191, 1, 7, 242, 2, 5, 
/* out0015_had-eta15-phi0*/	9, 1, 3, 5, 1, 8, 16, 1, 9, 16, 1, 10, 12, 3, 4, 16, 3, 7, 4, 190, 2, 7, 242, 1, 4, 242, 2, 1, 
/* out0016_had-eta16-phi0*/	7, 1, 2, 11, 1, 3, 2, 1, 6, 1, 1, 10, 4, 190, 1, 4, 190, 2, 3, 242, 1, 1, 
/* out0017_had-eta17-phi0*/	6, 1, 1, 3, 1, 2, 5, 1, 6, 15, 1, 7, 5, 190, 1, 5, 241, 1, 2, 
/* out0018_had-eta18-phi0*/	6, 0, 3, 16, 0, 4, 2, 1, 4, 16, 1, 7, 10, 190, 1, 1, 241, 1, 1, 
/* out0019_had-eta19-phi0*/	4, 0, 1, 16, 0, 2, 1, 0, 4, 12, 0, 5, 16, 
/* out0020_had-eta0-phi1*/	1, 253, 0, 1, 
/* out0021_had-eta1-phi1*/	1, 253, 0, 5, 
/* out0022_had-eta2-phi1*/	7, 39, 0, 10, 39, 2, 2, 51, 2, 3, 52, 0, 3, 52, 1, 15, 252, 0, 2, 253, 0, 2, 
/* out0023_had-eta3-phi1*/	8, 38, 0, 8, 38, 2, 5, 39, 0, 6, 39, 1, 4, 50, 2, 1, 51, 1, 12, 51, 2, 11, 252, 0, 4, 
/* out0024_had-eta4-phi1*/	8, 37, 0, 5, 37, 2, 5, 38, 0, 8, 38, 1, 6, 50, 1, 6, 50, 2, 8, 251, 0, 3, 252, 0, 2, 
/* out0025_had-eta5-phi1*/	8, 36, 0, 1, 36, 2, 3, 37, 0, 11, 37, 1, 8, 37, 2, 2, 49, 1, 2, 49, 2, 4, 251, 0, 4, 
/* out0026_had-eta6-phi1*/	6, 36, 0, 13, 36, 1, 6, 36, 2, 6, 49, 1, 1, 250, 0, 2, 251, 0, 1, 
/* out0027_had-eta7-phi1*/	5, 35, 0, 4, 35, 2, 11, 36, 0, 1, 36, 1, 5, 250, 0, 3, 
/* out0028_had-eta8-phi1*/	9, 34, 2, 1, 35, 0, 3, 35, 1, 13, 35, 2, 1, 189, 1, 9, 193, 0, 1, 239, 2, 1, 245, 0, 8, 250, 0, 2, 
/* out0029_had-eta9-phi1*/	13, 34, 0, 1, 34, 1, 1, 34, 2, 13, 188, 2, 7, 189, 1, 4, 193, 0, 7, 239, 1, 3, 239, 2, 4, 244, 0, 2, 244, 2, 3, 245, 0, 8, 245, 1, 4, 250, 0, 1, 
/* out0030_had-eta10-phi1*/	12, 9, 8, 1, 24, 0, 1, 34, 1, 11, 188, 1, 7, 188, 2, 3, 192, 0, 4, 192, 2, 1, 193, 0, 1, 193, 1, 3, 244, 0, 12, 244, 1, 2, 244, 2, 2, 
/* out0031_had-eta11-phi1*/	14, 9, 8, 15, 9, 9, 3, 9, 10, 7, 9, 11, 10, 24, 0, 1, 187, 2, 4, 188, 1, 1, 192, 0, 8, 192, 1, 2, 237, 2, 1, 243, 0, 2, 243, 2, 5, 244, 0, 1, 244, 1, 4, 
/* out0032_had-eta12-phi1*/	15, 3, 0, 1, 3, 3, 1, 9, 4, 5, 9, 5, 14, 9, 6, 7, 9, 10, 2, 9, 11, 3, 187, 1, 3, 187, 2, 2, 191, 0, 3, 191, 2, 2, 192, 1, 1, 243, 0, 6, 243, 1, 3, 243, 2, 3, 
/* out0033_had-eta13-phi1*/	10, 3, 0, 13, 3, 1, 1, 8, 8, 7, 9, 4, 7, 191, 0, 9, 191, 1, 2, 191, 2, 2, 242, 2, 3, 243, 0, 1, 243, 1, 6, 
/* out0034_had-eta14-phi1*/	11, 3, 0, 1, 3, 1, 4, 8, 5, 1, 8, 8, 3, 8, 11, 15, 186, 2, 1, 190, 2, 1, 191, 0, 3, 191, 1, 3, 242, 0, 1, 242, 2, 6, 
/* out0035_had-eta15-phi1*/	8, 1, 0, 1, 1, 3, 6, 8, 4, 2, 8, 5, 12, 190, 0, 4, 190, 2, 3, 242, 0, 1, 242, 1, 6, 
/* out0036_had-eta16-phi1*/	9, 1, 0, 11, 1, 1, 1, 1, 3, 3, 8, 4, 1, 190, 0, 5, 190, 1, 1, 190, 2, 1, 241, 1, 3, 242, 1, 3, 
/* out0037_had-eta17-phi1*/	7, 1, 0, 3, 1, 1, 8, 2, 8, 1, 2, 11, 1, 190, 0, 1, 190, 1, 4, 241, 1, 5, 
/* out0038_had-eta18-phi1*/	7, 0, 2, 5, 0, 4, 1, 1, 1, 4, 1, 7, 1, 2, 5, 2, 2, 11, 4, 241, 1, 1, 
/* out0039_had-eta19-phi1*/	3, 0, 2, 9, 0, 4, 1, 2, 5, 1, 
/* out0040_had-eta0-phi2*/	1, 257, 0, 1, 
/* out0041_had-eta1-phi2*/	1, 257, 0, 5, 
/* out0042_had-eta2-phi2*/	9, 51, 0, 1, 51, 2, 1, 52, 0, 13, 52, 1, 1, 91, 0, 5, 91, 1, 9, 91, 2, 16, 256, 0, 2, 257, 0, 2, 
/* out0043_had-eta3-phi2*/	9, 50, 0, 1, 50, 2, 2, 51, 0, 15, 51, 1, 4, 51, 2, 1, 90, 1, 6, 90, 2, 12, 91, 1, 6, 256, 0, 4, 
/* out0044_had-eta4-phi2*/	8, 50, 0, 15, 50, 1, 9, 50, 2, 5, 89, 1, 1, 89, 2, 5, 90, 1, 3, 255, 0, 3, 256, 0, 2, 
/* out0045_had-eta5-phi2*/	6, 49, 0, 12, 49, 1, 5, 49, 2, 12, 50, 1, 1, 89, 1, 1, 255, 0, 4, 
/* out0046_had-eta6-phi2*/	7, 36, 0, 1, 48, 0, 2, 48, 2, 14, 49, 0, 1, 49, 1, 8, 254, 0, 2, 255, 0, 1, 
/* out0047_had-eta7-phi2*/	6, 35, 0, 4, 47, 2, 2, 48, 0, 1, 48, 1, 13, 48, 2, 2, 254, 0, 3, 
/* out0048_had-eta8-phi2*/	9, 35, 0, 5, 47, 1, 3, 47, 2, 9, 183, 2, 6, 189, 0, 15, 189, 1, 1, 239, 0, 2, 239, 2, 6, 254, 0, 2, 
/* out0049_had-eta9-phi2*/	13, 34, 0, 10, 46, 2, 1, 47, 1, 4, 183, 1, 3, 183, 2, 2, 188, 0, 7, 188, 2, 5, 189, 0, 1, 189, 1, 2, 239, 0, 6, 239, 1, 8, 239, 2, 5, 254, 0, 1, 
/* out0050_had-eta10-phi2*/	12, 9, 3, 1, 9, 9, 4, 34, 0, 5, 34, 1, 3, 46, 1, 1, 46, 2, 2, 188, 0, 7, 188, 1, 7, 188, 2, 1, 237, 2, 11, 239, 1, 4, 244, 0, 1, 
/* out0051_had-eta11-phi2*/	11, 9, 0, 1, 9, 2, 9, 9, 3, 15, 9, 9, 9, 9, 10, 6, 187, 0, 3, 187, 2, 9, 188, 1, 1, 237, 1, 9, 237, 2, 3, 243, 0, 1, 
/* out0052_had-eta12-phi2*/	12, 9, 1, 7, 9, 2, 7, 9, 4, 1, 9, 6, 9, 9, 7, 10, 9, 10, 1, 187, 0, 1, 187, 1, 8, 187, 2, 1, 236, 2, 4, 237, 1, 2, 243, 0, 5, 
/* out0053_had-eta13-phi2*/	11, 8, 8, 6, 8, 9, 13, 8, 10, 1, 9, 4, 3, 9, 7, 5, 186, 2, 6, 187, 1, 3, 236, 1, 3, 236, 2, 3, 242, 0, 1, 243, 0, 1, 
/* out0054_had-eta14-phi2*/	9, 8, 2, 3, 8, 6, 4, 8, 9, 1, 8, 10, 15, 8, 11, 1, 186, 1, 3, 186, 2, 5, 236, 1, 1, 242, 0, 7, 
/* out0055_had-eta15-phi2*/	8, 8, 4, 4, 8, 5, 3, 8, 6, 9, 8, 7, 3, 186, 1, 5, 190, 0, 2, 242, 0, 5, 242, 1, 1, 
/* out0056_had-eta16-phi2*/	8, 1, 0, 1, 2, 8, 7, 8, 4, 8, 185, 2, 2, 190, 0, 3, 241, 0, 2, 241, 1, 2, 242, 1, 1, 
/* out0057_had-eta17-phi2*/	9, 2, 8, 7, 2, 10, 1, 2, 11, 6, 185, 1, 1, 185, 2, 2, 190, 0, 1, 190, 1, 1, 241, 0, 6, 241, 1, 2, 
/* out0058_had-eta18-phi2*/	4, 2, 5, 4, 2, 6, 1, 2, 10, 2, 2, 11, 5, 
/* out0059_had-eta19-phi2*/	4, 0, 0, 16, 0, 2, 1, 2, 4, 2, 2, 5, 7, 
/* out0060_had-eta0-phi3*/	1, 257, 0, 1, 
/* out0061_had-eta1-phi3*/	1, 257, 0, 5, 
/* out0062_had-eta2-phi3*/	7, 91, 0, 10, 102, 0, 4, 102, 1, 1, 102, 2, 15, 104, 2, 3, 256, 0, 2, 257, 0, 2, 
/* out0063_had-eta3-phi3*/	9, 90, 0, 16, 90, 1, 3, 90, 2, 4, 91, 0, 1, 91, 1, 1, 100, 2, 9, 102, 1, 13, 102, 2, 1, 256, 0, 4, 
/* out0064_had-eta4-phi3*/	8, 89, 0, 14, 89, 1, 4, 89, 2, 11, 90, 1, 4, 100, 1, 4, 100, 2, 1, 255, 0, 3, 256, 0, 2, 
/* out0065_had-eta5-phi3*/	6, 49, 0, 3, 88, 0, 3, 88, 2, 14, 89, 0, 1, 89, 1, 10, 255, 0, 4, 
/* out0066_had-eta6-phi3*/	6, 48, 0, 7, 87, 2, 2, 88, 1, 13, 88, 2, 2, 254, 0, 2, 255, 0, 1, 
/* out0067_had-eta7-phi3*/	7, 47, 0, 2, 47, 2, 2, 48, 0, 6, 48, 1, 3, 87, 1, 4, 87, 2, 6, 254, 0, 3, 
/* out0068_had-eta8-phi3*/	7, 47, 0, 11, 47, 1, 3, 47, 2, 3, 183, 0, 7, 183, 2, 8, 239, 0, 1, 254, 0, 2, 
/* out0069_had-eta9-phi3*/	10, 46, 2, 7, 47, 0, 1, 47, 1, 6, 182, 2, 3, 183, 0, 3, 183, 1, 13, 188, 0, 1, 239, 0, 7, 240, 2, 11, 254, 0, 1, 
/* out0070_had-eta10-phi3*/	10, 46, 0, 1, 46, 1, 5, 46, 2, 6, 182, 1, 3, 182, 2, 11, 188, 0, 1, 237, 0, 8, 237, 2, 1, 239, 1, 1, 240, 1, 6, 
/* out0071_had-eta11-phi3*/	9, 9, 0, 11, 10, 8, 7, 46, 1, 6, 181, 2, 1, 182, 1, 6, 187, 0, 6, 237, 0, 8, 237, 1, 4, 238, 2, 1, 
/* out0072_had-eta12-phi3*/	11, 9, 0, 4, 9, 1, 9, 10, 5, 1, 10, 8, 6, 10, 11, 15, 181, 2, 3, 187, 0, 6, 187, 1, 1, 236, 0, 3, 236, 2, 7, 237, 1, 1, 
/* out0073_had-eta13-phi3*/	13, 8, 0, 2, 8, 3, 12, 8, 9, 2, 9, 7, 1, 10, 4, 1, 10, 5, 10, 181, 1, 1, 186, 0, 4, 186, 2, 3, 187, 1, 1, 236, 0, 2, 236, 1, 6, 236, 2, 2, 
/* out0074_had-eta14-phi3*/	10, 8, 0, 5, 8, 1, 4, 8, 2, 11, 8, 3, 4, 186, 0, 5, 186, 1, 2, 186, 2, 1, 235, 2, 3, 236, 1, 4, 242, 0, 1, 
/* out0075_had-eta15-phi3*/	7, 8, 1, 7, 8, 2, 2, 8, 6, 3, 8, 7, 9, 185, 2, 1, 186, 1, 5, 235, 2, 6, 
/* out0076_had-eta16-phi3*/	7, 2, 8, 1, 2, 9, 11, 8, 4, 1, 8, 7, 4, 185, 2, 5, 235, 1, 4, 241, 0, 2, 
/* out0077_had-eta17-phi3*/	7, 2, 2, 1, 2, 9, 3, 2, 10, 10, 185, 1, 4, 185, 2, 3, 235, 1, 1, 241, 0, 6, 
/* out0078_had-eta18-phi3*/	4, 2, 2, 1, 2, 6, 8, 2, 10, 3, 185, 1, 2, 
/* out0079_had-eta19-phi3*/	4, 2, 4, 4, 2, 5, 2, 2, 6, 3, 2, 7, 2, 
/* out0080_had-eta0-phi4*/	1, 261, 0, 1, 
/* out0081_had-eta1-phi4*/	1, 261, 0, 5, 
/* out0082_had-eta2-phi4*/	8, 102, 0, 9, 103, 0, 2, 103, 2, 11, 104, 0, 16, 104, 1, 16, 104, 2, 13, 260, 0, 2, 261, 0, 2, 
/* out0083_had-eta3-phi4*/	10, 100, 0, 13, 100, 1, 1, 100, 2, 6, 101, 2, 3, 102, 0, 3, 102, 1, 2, 103, 0, 1, 103, 1, 11, 103, 2, 5, 260, 0, 4, 
/* out0084_had-eta4-phi4*/	9, 89, 0, 1, 99, 0, 7, 99, 2, 13, 100, 0, 3, 100, 1, 11, 101, 1, 1, 101, 2, 2, 259, 0, 3, 260, 0, 2, 
/* out0085_had-eta5-phi4*/	6, 88, 0, 8, 98, 2, 5, 99, 0, 1, 99, 1, 14, 99, 2, 3, 259, 0, 4, 
/* out0086_had-eta6-phi4*/	8, 87, 0, 4, 87, 2, 4, 88, 0, 5, 88, 1, 3, 98, 1, 4, 98, 2, 5, 258, 0, 2, 259, 0, 1, 
/* out0087_had-eta7-phi4*/	4, 87, 0, 9, 87, 1, 9, 87, 2, 4, 258, 0, 3, 
/* out0088_had-eta8-phi4*/	8, 47, 0, 2, 86, 2, 13, 87, 1, 3, 183, 0, 3, 184, 2, 6, 240, 0, 1, 240, 2, 1, 258, 0, 2, 
/* out0089_had-eta9-phi4*/	12, 46, 0, 5, 86, 1, 8, 86, 2, 2, 182, 0, 2, 182, 2, 1, 183, 0, 3, 184, 1, 6, 184, 2, 8, 240, 0, 12, 240, 1, 1, 240, 2, 4, 258, 0, 1, 
/* out0090_had-eta10-phi4*/	9, 46, 0, 10, 46, 1, 1, 139, 2, 1, 182, 0, 13, 182, 1, 2, 182, 2, 1, 238, 2, 6, 240, 0, 2, 240, 1, 9, 
/* out0091_had-eta11-phi4*/	11, 10, 3, 6, 10, 8, 3, 10, 9, 15, 10, 10, 1, 46, 1, 3, 181, 0, 1, 181, 2, 6, 182, 0, 1, 182, 1, 5, 238, 1, 4, 238, 2, 9, 
/* out0092_had-eta12-phi4*/	11, 10, 2, 8, 10, 6, 8, 10, 9, 1, 10, 10, 15, 10, 11, 1, 181, 0, 1, 181, 1, 3, 181, 2, 6, 236, 0, 5, 238, 1, 6, 246, 2, 1, 
/* out0093_had-eta13-phi4*/	9, 10, 4, 13, 10, 5, 5, 10, 6, 6, 10, 7, 3, 181, 1, 7, 186, 0, 2, 236, 0, 6, 236, 1, 1, 246, 2, 2, 
/* out0094_had-eta14-phi4*/	9, 8, 0, 9, 10, 4, 1, 14, 8, 10, 14, 11, 1, 175, 2, 3, 186, 0, 4, 235, 0, 2, 235, 2, 4, 236, 1, 1, 
/* out0095_had-eta15-phi4*/	12, 8, 1, 5, 14, 5, 2, 14, 11, 11, 175, 1, 1, 175, 2, 1, 185, 0, 1, 185, 2, 1, 186, 0, 1, 186, 1, 1, 235, 0, 3, 235, 1, 1, 235, 2, 3, 
/* out0096_had-eta16-phi4*/	6, 2, 3, 10, 2, 9, 2, 14, 5, 4, 185, 0, 4, 185, 2, 2, 235, 1, 5, 
/* out0097_had-eta17-phi4*/	5, 2, 2, 7, 2, 3, 6, 185, 0, 2, 185, 1, 3, 235, 1, 2, 
/* out0098_had-eta18-phi4*/	4, 2, 1, 2, 2, 2, 7, 2, 6, 3, 185, 1, 4, 
/* out0099_had-eta19-phi4*/	3, 2, 4, 10, 2, 6, 1, 2, 7, 9, 
/* out0100_had-eta0-phi5*/	1, 261, 0, 1, 
/* out0101_had-eta1-phi5*/	1, 261, 0, 5, 
/* out0102_had-eta2-phi5*/	4, 103, 0, 7, 114, 2, 6, 260, 0, 2, 261, 0, 2, 
/* out0103_had-eta3-phi5*/	7, 101, 0, 11, 101, 2, 9, 103, 0, 6, 103, 1, 5, 114, 1, 8, 114, 2, 10, 260, 0, 4, 
/* out0104_had-eta4-phi5*/	7, 99, 0, 5, 101, 0, 5, 101, 1, 15, 101, 2, 2, 112, 2, 11, 259, 0, 3, 260, 0, 2, 
/* out0105_had-eta5-phi5*/	7, 98, 0, 8, 98, 2, 4, 99, 0, 3, 99, 1, 2, 112, 1, 8, 112, 2, 5, 259, 0, 4, 
/* out0106_had-eta6-phi5*/	6, 98, 0, 8, 98, 1, 12, 98, 2, 2, 122, 2, 4, 258, 0, 2, 259, 0, 1, 
/* out0107_had-eta7-phi5*/	4, 87, 0, 3, 122, 1, 5, 122, 2, 12, 258, 0, 3, 
/* out0108_had-eta8-phi5*/	6, 86, 0, 13, 86, 2, 1, 122, 1, 3, 184, 0, 6, 184, 2, 1, 258, 0, 2, 
/* out0109_had-eta9-phi5*/	10, 86, 0, 3, 86, 1, 8, 139, 2, 3, 177, 2, 1, 184, 0, 10, 184, 1, 9, 184, 2, 1, 240, 0, 1, 248, 2, 13, 258, 0, 1, 
/* out0110_had-eta10-phi5*/	7, 139, 1, 1, 139, 2, 11, 177, 2, 13, 184, 1, 1, 238, 0, 5, 248, 1, 8, 248, 2, 3, 
/* out0111_had-eta11-phi5*/	9, 10, 0, 5, 10, 3, 8, 139, 1, 6, 139, 2, 1, 177, 1, 7, 177, 2, 1, 181, 0, 4, 238, 0, 11, 238, 1, 2, 
/* out0112_had-eta12-phi5*/	9, 10, 0, 11, 10, 1, 11, 10, 2, 8, 10, 3, 2, 10, 6, 1, 181, 0, 9, 181, 1, 1, 238, 1, 4, 246, 2, 6, 
/* out0113_had-eta13-phi5*/	11, 10, 1, 5, 10, 4, 1, 10, 6, 1, 10, 7, 13, 14, 8, 1, 14, 9, 6, 175, 2, 4, 181, 0, 1, 181, 1, 4, 246, 1, 2, 246, 2, 7, 
/* out0114_had-eta14-phi5*/	7, 14, 8, 5, 14, 9, 9, 14, 10, 8, 14, 11, 1, 175, 2, 7, 235, 0, 3, 246, 1, 5, 
/* out0115_had-eta15-phi5*/	7, 14, 5, 3, 14, 6, 7, 14, 10, 7, 14, 11, 3, 175, 1, 6, 175, 2, 1, 235, 0, 6, 
/* out0116_had-eta16-phi5*/	7, 2, 0, 2, 14, 4, 7, 14, 5, 7, 175, 1, 1, 185, 0, 4, 235, 0, 2, 235, 1, 3, 
/* out0117_had-eta17-phi5*/	3, 2, 0, 12, 2, 1, 1, 185, 0, 4, 
/* out0118_had-eta18-phi5*/	4, 2, 0, 2, 2, 1, 9, 185, 0, 1, 185, 1, 2, 
/* out0119_had-eta19-phi5*/	2, 2, 1, 4, 2, 7, 5, 
/* out0120_had-eta0-phi6*/	1, 265, 0, 1, 
/* out0121_had-eta1-phi6*/	1, 265, 0, 5, 
/* out0122_had-eta2-phi6*/	4, 114, 0, 6, 115, 2, 7, 264, 0, 2, 265, 0, 2, 
/* out0123_had-eta3-phi6*/	7, 113, 0, 9, 113, 2, 11, 114, 0, 10, 114, 1, 8, 115, 1, 4, 115, 2, 6, 264, 0, 4, 
/* out0124_had-eta4-phi6*/	7, 112, 0, 11, 113, 0, 2, 113, 1, 15, 113, 2, 5, 124, 2, 5, 263, 0, 3, 264, 0, 2, 
/* out0125_had-eta5-phi6*/	7, 112, 0, 5, 112, 1, 8, 123, 0, 4, 123, 2, 8, 124, 1, 2, 124, 2, 3, 263, 0, 4, 
/* out0126_had-eta6-phi6*/	6, 122, 0, 4, 123, 0, 2, 123, 1, 12, 123, 2, 8, 262, 0, 2, 263, 0, 1, 
/* out0127_had-eta7-phi6*/	4, 122, 0, 12, 122, 1, 5, 141, 2, 3, 262, 0, 3, 
/* out0128_had-eta8-phi6*/	6, 122, 1, 3, 140, 0, 1, 140, 2, 13, 179, 0, 1, 179, 2, 6, 262, 0, 2, 
/* out0129_had-eta9-phi6*/	10, 139, 0, 4, 140, 1, 8, 140, 2, 3, 177, 0, 1, 179, 0, 1, 179, 1, 9, 179, 2, 10, 248, 0, 13, 249, 2, 1, 262, 0, 1, 
/* out0130_had-eta10-phi6*/	9, 139, 0, 11, 139, 1, 2, 177, 0, 14, 177, 1, 1, 177, 2, 1, 179, 1, 1, 247, 2, 5, 248, 0, 3, 248, 1, 8, 
/* out0131_had-eta11-phi6*/	8, 15, 8, 5, 15, 9, 8, 139, 1, 7, 176, 2, 4, 177, 0, 1, 177, 1, 8, 247, 1, 2, 247, 2, 11, 
/* out0132_had-eta12-phi6*/	9, 15, 6, 1, 15, 8, 11, 15, 9, 2, 15, 10, 8, 15, 11, 11, 176, 1, 1, 176, 2, 9, 246, 0, 6, 247, 1, 4, 
/* out0133_had-eta13-phi6*/	12, 14, 0, 1, 14, 3, 7, 14, 9, 1, 15, 4, 1, 15, 5, 13, 15, 6, 1, 15, 11, 5, 175, 0, 4, 176, 1, 4, 176, 2, 1, 246, 0, 7, 246, 1, 3, 
/* out0134_had-eta14-phi6*/	8, 14, 0, 3, 14, 1, 1, 14, 2, 9, 14, 3, 9, 14, 10, 1, 175, 0, 7, 231, 2, 3, 246, 1, 5, 
/* out0135_had-eta15-phi6*/	7, 14, 1, 2, 14, 2, 7, 14, 6, 8, 14, 7, 3, 175, 0, 1, 175, 1, 6, 231, 2, 6, 
/* out0136_had-eta16-phi6*/	8, 14, 4, 8, 14, 6, 1, 14, 7, 6, 18, 8, 2, 170, 2, 4, 175, 1, 1, 231, 1, 3, 231, 2, 2, 
/* out0137_had-eta17-phi6*/	4, 14, 4, 1, 18, 8, 12, 18, 11, 1, 170, 2, 4, 
/* out0138_had-eta18-phi6*/	4, 18, 8, 2, 18, 11, 9, 170, 1, 2, 170, 2, 1, 
/* out0139_had-eta19-phi6*/	2, 18, 5, 5, 18, 11, 4, 
/* out0140_had-eta0-phi7*/	1, 265, 0, 1, 
/* out0141_had-eta1-phi7*/	1, 265, 0, 5, 
/* out0142_had-eta2-phi7*/	8, 115, 0, 11, 115, 2, 2, 116, 0, 13, 116, 1, 16, 116, 2, 16, 126, 2, 9, 264, 0, 2, 265, 0, 2, 
/* out0143_had-eta3-phi7*/	10, 113, 0, 3, 115, 0, 5, 115, 1, 12, 115, 2, 1, 125, 0, 6, 125, 1, 1, 125, 2, 13, 126, 1, 2, 126, 2, 3, 264, 0, 4, 
/* out0144_had-eta4-phi7*/	9, 113, 0, 2, 113, 1, 1, 124, 0, 13, 124, 2, 7, 125, 1, 11, 125, 2, 3, 143, 2, 1, 263, 0, 3, 264, 0, 2, 
/* out0145_had-eta5-phi7*/	6, 123, 0, 5, 124, 0, 3, 124, 1, 14, 124, 2, 1, 142, 2, 8, 263, 0, 4, 
/* out0146_had-eta6-phi7*/	8, 123, 0, 5, 123, 1, 4, 141, 0, 4, 141, 2, 4, 142, 1, 3, 142, 2, 5, 262, 0, 2, 263, 0, 1, 
/* out0147_had-eta7-phi7*/	4, 141, 0, 4, 141, 1, 9, 141, 2, 9, 262, 0, 3, 
/* out0148_had-eta8-phi7*/	8, 61, 2, 2, 140, 0, 13, 141, 1, 3, 179, 0, 6, 180, 2, 3, 249, 0, 1, 249, 2, 1, 262, 0, 2, 
/* out0149_had-eta9-phi7*/	12, 60, 2, 5, 140, 0, 2, 140, 1, 8, 178, 0, 1, 178, 2, 2, 179, 0, 8, 179, 1, 6, 180, 2, 3, 249, 0, 4, 249, 1, 1, 249, 2, 12, 262, 0, 1, 
/* out0150_had-eta10-phi7*/	9, 60, 1, 1, 60, 2, 10, 139, 0, 1, 178, 0, 1, 178, 1, 2, 178, 2, 13, 247, 0, 6, 249, 1, 9, 249, 2, 2, 
/* out0151_had-eta11-phi7*/	11, 15, 0, 3, 15, 2, 1, 15, 3, 15, 15, 9, 6, 60, 1, 3, 176, 0, 6, 176, 2, 1, 178, 1, 5, 178, 2, 1, 247, 0, 9, 247, 1, 4, 
/* out0152_had-eta12-phi7*/	11, 15, 1, 1, 15, 2, 15, 15, 3, 1, 15, 6, 8, 15, 10, 8, 176, 0, 6, 176, 1, 3, 176, 2, 1, 232, 2, 5, 246, 0, 1, 247, 1, 6, 
/* out0153_had-eta13-phi7*/	9, 15, 4, 13, 15, 5, 3, 15, 6, 6, 15, 7, 5, 171, 2, 2, 176, 1, 7, 232, 1, 1, 232, 2, 6, 246, 0, 2, 
/* out0154_had-eta14-phi7*/	10, 14, 0, 12, 14, 1, 1, 15, 4, 1, 19, 8, 9, 171, 2, 4, 175, 0, 3, 231, 0, 4, 231, 2, 2, 232, 1, 1, 246, 1, 1, 
/* out0155_had-eta15-phi7*/	12, 14, 1, 12, 14, 7, 2, 19, 11, 5, 170, 0, 1, 170, 2, 1, 171, 1, 1, 171, 2, 1, 175, 0, 1, 175, 1, 1, 231, 0, 3, 231, 1, 1, 231, 2, 3, 
/* out0156_had-eta16-phi7*/	6, 14, 7, 5, 18, 3, 2, 18, 9, 10, 170, 0, 2, 170, 2, 4, 231, 1, 5, 
/* out0157_had-eta17-phi7*/	5, 18, 9, 6, 18, 10, 7, 170, 1, 3, 170, 2, 2, 231, 1, 2, 
/* out0158_had-eta18-phi7*/	4, 18, 6, 3, 18, 10, 7, 18, 11, 2, 170, 1, 4, 
/* out0159_had-eta19-phi7*/	3, 18, 4, 10, 18, 5, 9, 18, 6, 1, 
/* out0160_had-eta0-phi8*/	1, 269, 0, 1, 
/* out0161_had-eta1-phi8*/	1, 269, 0, 5, 
/* out0162_had-eta2-phi8*/	7, 116, 0, 3, 126, 0, 15, 126, 1, 1, 126, 2, 4, 145, 2, 10, 268, 0, 2, 269, 0, 2, 
/* out0163_had-eta3-phi8*/	9, 125, 0, 9, 126, 0, 1, 126, 1, 13, 144, 0, 4, 144, 1, 3, 144, 2, 16, 145, 1, 1, 145, 2, 1, 268, 0, 4, 
/* out0164_had-eta4-phi8*/	8, 125, 0, 1, 125, 1, 4, 143, 0, 11, 143, 1, 4, 143, 2, 14, 144, 1, 4, 267, 0, 3, 268, 0, 2, 
/* out0165_had-eta5-phi8*/	6, 63, 2, 3, 142, 0, 14, 142, 2, 3, 143, 1, 10, 143, 2, 1, 267, 0, 4, 
/* out0166_had-eta6-phi8*/	6, 62, 2, 7, 141, 0, 2, 142, 0, 2, 142, 1, 13, 266, 0, 2, 267, 0, 1, 
/* out0167_had-eta7-phi8*/	7, 61, 0, 2, 61, 2, 2, 62, 1, 3, 62, 2, 6, 141, 0, 6, 141, 1, 4, 266, 0, 3, 
/* out0168_had-eta8-phi8*/	7, 61, 0, 3, 61, 1, 3, 61, 2, 11, 180, 0, 8, 180, 2, 7, 234, 2, 1, 266, 0, 2, 
/* out0169_had-eta9-phi8*/	10, 60, 0, 7, 61, 1, 6, 61, 2, 1, 173, 2, 1, 178, 0, 3, 180, 1, 13, 180, 2, 3, 234, 2, 7, 249, 0, 11, 266, 0, 1, 
/* out0170_had-eta10-phi8*/	10, 60, 0, 6, 60, 1, 5, 60, 2, 1, 173, 2, 1, 178, 0, 11, 178, 1, 3, 233, 0, 1, 233, 2, 8, 234, 1, 1, 249, 1, 6, 
/* out0171_had-eta11-phi8*/	9, 15, 0, 7, 20, 8, 11, 60, 1, 6, 172, 2, 6, 176, 0, 1, 178, 1, 6, 233, 1, 4, 233, 2, 8, 247, 0, 1, 
/* out0172_had-eta12-phi8*/	11, 15, 0, 6, 15, 1, 15, 15, 7, 1, 20, 8, 4, 20, 11, 9, 172, 1, 1, 172, 2, 6, 176, 0, 3, 232, 0, 7, 232, 2, 3, 233, 1, 1, 
/* out0173_had-eta13-phi8*/	13, 15, 4, 1, 15, 7, 10, 19, 3, 2, 19, 8, 2, 19, 9, 12, 20, 5, 1, 171, 0, 3, 171, 2, 4, 172, 1, 1, 176, 1, 1, 232, 0, 2, 232, 1, 6, 232, 2, 2, 
/* out0174_had-eta14-phi8*/	10, 19, 8, 5, 19, 9, 4, 19, 10, 11, 19, 11, 4, 171, 0, 1, 171, 1, 2, 171, 2, 5, 227, 2, 1, 231, 0, 3, 232, 1, 4, 
/* out0175_had-eta15-phi8*/	7, 19, 5, 9, 19, 6, 3, 19, 10, 2, 19, 11, 7, 170, 0, 1, 171, 1, 5, 231, 0, 6, 
/* out0176_had-eta16-phi8*/	7, 18, 0, 1, 18, 3, 11, 19, 4, 1, 19, 5, 4, 170, 0, 5, 226, 1, 2, 231, 1, 4, 
/* out0177_had-eta17-phi8*/	7, 18, 2, 10, 18, 3, 3, 18, 10, 1, 170, 0, 3, 170, 1, 4, 226, 1, 6, 231, 1, 1, 
/* out0178_had-eta18-phi8*/	4, 18, 2, 3, 18, 6, 8, 18, 10, 1, 170, 1, 2, 
/* out0179_had-eta19-phi8*/	4, 18, 4, 4, 18, 5, 2, 18, 6, 3, 18, 7, 2, 
/* out0180_had-eta0-phi9*/	1, 269, 0, 1, 
/* out0181_had-eta1-phi9*/	1, 269, 0, 5, 
/* out0182_had-eta2-phi9*/	9, 65, 0, 1, 65, 2, 1, 66, 0, 1, 66, 1, 13, 145, 0, 16, 145, 1, 9, 145, 2, 5, 268, 0, 2, 269, 0, 2, 
/* out0183_had-eta3-phi9*/	9, 64, 0, 2, 64, 2, 1, 65, 0, 1, 65, 1, 4, 65, 2, 15, 144, 0, 12, 144, 1, 6, 145, 1, 6, 268, 0, 4, 
/* out0184_had-eta4-phi9*/	8, 64, 0, 5, 64, 1, 9, 64, 2, 15, 143, 0, 5, 143, 1, 1, 144, 1, 3, 267, 0, 3, 268, 0, 2, 
/* out0185_had-eta5-phi9*/	6, 63, 0, 12, 63, 1, 5, 63, 2, 12, 64, 1, 1, 143, 1, 1, 267, 0, 4, 
/* out0186_had-eta6-phi9*/	7, 62, 0, 14, 62, 2, 2, 63, 1, 8, 63, 2, 1, 76, 2, 1, 266, 0, 2, 267, 0, 1, 
/* out0187_had-eta7-phi9*/	6, 61, 0, 2, 62, 0, 2, 62, 1, 13, 62, 2, 1, 75, 2, 4, 266, 0, 3, 
/* out0188_had-eta8-phi9*/	9, 61, 0, 9, 61, 1, 3, 75, 2, 5, 174, 0, 1, 174, 1, 15, 180, 0, 6, 234, 0, 6, 234, 2, 2, 266, 0, 2, 
/* out0189_had-eta9-phi9*/	13, 60, 0, 1, 61, 1, 4, 74, 2, 10, 173, 0, 5, 173, 2, 7, 174, 0, 2, 174, 1, 1, 180, 0, 2, 180, 1, 3, 234, 0, 5, 234, 1, 8, 234, 2, 6, 266, 0, 1, 
/* out0190_had-eta10-phi9*/	12, 20, 3, 4, 20, 9, 1, 60, 0, 2, 60, 1, 1, 74, 1, 3, 74, 2, 5, 173, 0, 1, 173, 1, 7, 173, 2, 7, 229, 2, 1, 233, 0, 11, 234, 1, 4, 
/* out0191_had-eta11-phi9*/	11, 20, 2, 6, 20, 3, 9, 20, 8, 1, 20, 9, 15, 20, 10, 9, 172, 0, 9, 172, 2, 3, 173, 1, 1, 228, 2, 1, 233, 0, 3, 233, 1, 9, 
/* out0192_had-eta12-phi9*/	12, 20, 2, 1, 20, 4, 1, 20, 5, 10, 20, 6, 9, 20, 10, 7, 20, 11, 7, 172, 0, 1, 172, 1, 8, 172, 2, 1, 228, 2, 5, 232, 0, 4, 233, 1, 2, 
/* out0193_had-eta13-phi9*/	11, 19, 0, 6, 19, 2, 1, 19, 3, 13, 20, 4, 3, 20, 5, 5, 171, 0, 6, 172, 1, 3, 227, 2, 1, 228, 2, 1, 232, 0, 3, 232, 1, 3, 
/* out0194_had-eta14-phi9*/	9, 19, 1, 1, 19, 2, 15, 19, 3, 1, 19, 6, 4, 19, 10, 3, 171, 0, 5, 171, 1, 3, 227, 2, 7, 232, 1, 1, 
/* out0195_had-eta15-phi9*/	8, 19, 4, 4, 19, 5, 3, 19, 6, 9, 19, 7, 3, 166, 2, 2, 171, 1, 5, 227, 1, 1, 227, 2, 5, 
/* out0196_had-eta16-phi9*/	7, 18, 0, 7, 19, 4, 8, 166, 2, 3, 170, 0, 2, 226, 0, 2, 226, 1, 2, 227, 1, 1, 
/* out0197_had-eta17-phi9*/	8, 18, 0, 7, 18, 1, 6, 18, 2, 1, 166, 2, 1, 170, 0, 2, 170, 1, 1, 226, 0, 2, 226, 1, 6, 
/* out0198_had-eta18-phi9*/	4, 18, 1, 5, 18, 2, 2, 18, 6, 1, 18, 7, 4, 
/* out0199_had-eta19-phi9*/	4, 4, 4, 16, 4, 5, 1, 18, 4, 2, 18, 7, 7, 
/* out0200_had-eta0-phi10*/	1, 273, 0, 1, 
/* out0201_had-eta1-phi10*/	1, 273, 0, 5, 
/* out0202_had-eta2-phi10*/	7, 65, 0, 3, 66, 0, 15, 66, 1, 3, 79, 0, 2, 79, 2, 10, 272, 0, 2, 273, 0, 2, 
/* out0203_had-eta3-phi10*/	8, 64, 0, 1, 65, 0, 11, 65, 1, 12, 78, 0, 5, 78, 2, 8, 79, 1, 4, 79, 2, 6, 272, 0, 4, 
/* out0204_had-eta4-phi10*/	8, 64, 0, 8, 64, 1, 6, 77, 0, 5, 77, 2, 5, 78, 1, 6, 78, 2, 8, 271, 0, 3, 272, 0, 2, 
/* out0205_had-eta5-phi10*/	8, 63, 0, 4, 63, 1, 2, 76, 0, 3, 76, 2, 1, 77, 0, 2, 77, 1, 8, 77, 2, 11, 271, 0, 4, 
/* out0206_had-eta6-phi10*/	6, 63, 1, 1, 76, 0, 6, 76, 1, 6, 76, 2, 13, 270, 0, 2, 271, 0, 1, 
/* out0207_had-eta7-phi10*/	5, 75, 0, 11, 75, 2, 4, 76, 1, 5, 76, 2, 1, 270, 0, 3, 
/* out0208_had-eta8-phi10*/	9, 74, 0, 1, 75, 0, 1, 75, 1, 13, 75, 2, 3, 169, 2, 1, 174, 0, 9, 230, 1, 8, 234, 0, 1, 270, 0, 2, 
/* out0209_had-eta9-phi10*/	13, 74, 0, 13, 74, 1, 1, 74, 2, 1, 169, 2, 7, 173, 0, 7, 174, 0, 4, 229, 0, 3, 229, 2, 2, 230, 0, 4, 230, 1, 8, 234, 0, 4, 234, 1, 3, 270, 0, 1, 
/* out0210_had-eta10-phi10*/	10, 20, 0, 1, 29, 2, 1, 74, 1, 11, 168, 2, 4, 169, 2, 1, 173, 0, 3, 173, 1, 7, 229, 0, 2, 229, 1, 2, 229, 2, 12, 
/* out0211_had-eta11-phi10*/	13, 20, 0, 15, 20, 1, 10, 20, 2, 7, 20, 3, 3, 29, 2, 1, 168, 2, 8, 172, 0, 4, 173, 1, 1, 228, 0, 5, 228, 2, 2, 229, 1, 4, 229, 2, 1, 233, 0, 1, 
/* out0212_had-eta12-phi10*/	14, 7, 9, 1, 20, 1, 3, 20, 2, 2, 20, 4, 5, 20, 6, 7, 20, 7, 14, 167, 0, 1, 167, 2, 3, 168, 1, 1, 172, 0, 2, 172, 1, 3, 228, 0, 3, 228, 1, 3, 228, 2, 6, 
/* out0213_had-eta13-phi10*/	7, 7, 8, 13, 19, 0, 7, 20, 4, 7, 167, 2, 9, 227, 0, 3, 228, 1, 6, 228, 2, 1, 
/* out0214_had-eta14-phi10*/	11, 7, 8, 1, 7, 11, 3, 19, 0, 3, 19, 1, 15, 19, 7, 1, 166, 0, 1, 167, 1, 2, 167, 2, 3, 171, 0, 1, 227, 0, 6, 227, 2, 1, 
/* out0215_had-eta15-phi10*/	8, 6, 8, 1, 6, 9, 4, 19, 4, 2, 19, 7, 12, 166, 0, 2, 166, 2, 4, 227, 1, 6, 227, 2, 1, 
/* out0216_had-eta16-phi10*/	8, 6, 8, 12, 6, 9, 3, 6, 11, 1, 19, 4, 1, 166, 1, 1, 166, 2, 5, 226, 0, 3, 227, 1, 3, 
/* out0217_had-eta17-phi10*/	7, 6, 8, 3, 6, 11, 7, 18, 0, 1, 18, 1, 1, 166, 1, 4, 166, 2, 1, 226, 0, 5, 
/* out0218_had-eta18-phi10*/	6, 4, 3, 1, 4, 5, 1, 6, 11, 3, 18, 1, 4, 18, 7, 2, 226, 0, 1, 
/* out0219_had-eta19-phi10*/	2, 4, 5, 9, 18, 7, 1, 
/* out0220_had-eta0-phi11*/	1, 273, 0, 1, 
/* out0221_had-eta1-phi11*/	1, 273, 0, 5, 
/* out0222_had-eta2-phi11*/	3, 79, 0, 14, 272, 0, 2, 273, 0, 2, 
/* out0223_had-eta3-phi11*/	3, 78, 0, 10, 79, 1, 12, 272, 0, 4, 
/* out0224_had-eta4-phi11*/	8, 33, 0, 4, 33, 1, 1, 33, 2, 15, 77, 0, 5, 78, 0, 1, 78, 1, 10, 271, 0, 3, 272, 0, 2, 
/* out0225_had-eta5-phi11*/	8, 32, 0, 4, 32, 2, 10, 33, 1, 3, 33, 2, 1, 76, 0, 1, 77, 0, 4, 77, 1, 8, 271, 0, 4, 
/* out0226_had-eta6-phi11*/	8, 31, 0, 3, 31, 2, 3, 32, 1, 4, 32, 2, 6, 76, 0, 6, 76, 1, 4, 270, 0, 2, 271, 0, 1, 
/* out0227_had-eta7-phi11*/	6, 31, 0, 1, 31, 1, 2, 31, 2, 13, 75, 0, 3, 76, 1, 1, 270, 0, 3, 
/* out0228_had-eta8-phi11*/	9, 30, 0, 4, 30, 2, 7, 31, 1, 1, 75, 0, 1, 75, 1, 3, 169, 0, 6, 169, 2, 1, 230, 0, 3, 270, 0, 2, 
/* out0229_had-eta9-phi11*/	10, 30, 1, 4, 30, 2, 9, 74, 0, 2, 169, 0, 6, 169, 1, 7, 169, 2, 6, 225, 2, 6, 229, 0, 4, 230, 0, 9, 270, 0, 1, 
/* out0230_had-eta10-phi11*/	10, 29, 0, 4, 29, 2, 7, 74, 1, 1, 168, 0, 9, 168, 2, 1, 169, 1, 5, 224, 2, 1, 225, 2, 1, 229, 0, 7, 229, 1, 6, 
/* out0231_had-eta11-phi11*/	9, 20, 1, 1, 29, 1, 2, 29, 2, 7, 168, 0, 3, 168, 1, 7, 168, 2, 3, 224, 2, 6, 228, 0, 3, 229, 1, 4, 
/* out0232_had-eta12-phi11*/	11, 7, 2, 1, 7, 3, 12, 7, 9, 10, 20, 1, 2, 20, 7, 2, 29, 1, 2, 167, 0, 7, 168, 1, 4, 224, 2, 1, 228, 0, 5, 228, 1, 4, 
/* out0233_had-eta13-phi11*/	12, 7, 2, 2, 7, 6, 1, 7, 8, 2, 7, 9, 5, 7, 10, 15, 7, 11, 3, 167, 0, 4, 167, 1, 3, 167, 2, 1, 223, 2, 5, 227, 0, 1, 228, 1, 3, 
/* out0234_had-eta14-phi11*/	8, 7, 5, 11, 7, 6, 2, 7, 10, 1, 7, 11, 10, 166, 0, 1, 167, 1, 7, 223, 2, 2, 227, 0, 5, 
/* out0235_had-eta15-phi11*/	8, 6, 2, 1, 6, 3, 12, 6, 9, 6, 7, 5, 1, 166, 0, 6, 222, 2, 2, 227, 0, 1, 227, 1, 4, 
/* out0236_had-eta16-phi11*/	7, 6, 2, 3, 6, 9, 3, 6, 10, 11, 166, 0, 2, 166, 1, 3, 222, 2, 4, 227, 1, 1, 
/* out0237_had-eta17-phi11*/	7, 6, 5, 2, 6, 6, 3, 6, 10, 5, 6, 11, 4, 166, 1, 4, 222, 2, 2, 226, 0, 2, 
/* out0238_had-eta18-phi11*/	4, 4, 3, 2, 6, 5, 9, 6, 11, 1, 226, 0, 1, 
/* out0239_had-eta19-phi11*/	4, 4, 2, 15, 4, 3, 9, 4, 5, 5, 4, 6, 16, 
/* out0240_had-eta0-phi12*/	1, 277, 0, 1, 
/* out0241_had-eta1-phi12*/	1, 277, 0, 5, 
/* out0242_had-eta2-phi12*/	4, 45, 0, 6, 45, 2, 8, 276, 0, 2, 277, 0, 2, 
/* out0243_had-eta3-phi12*/	5, 44, 0, 4, 44, 2, 7, 45, 1, 5, 45, 2, 8, 276, 0, 4, 
/* out0244_had-eta4-phi12*/	8, 33, 0, 12, 33, 1, 8, 43, 0, 2, 43, 2, 3, 44, 1, 2, 44, 2, 9, 275, 0, 3, 276, 0, 2, 
/* out0245_had-eta5-phi12*/	6, 32, 0, 12, 32, 1, 2, 33, 1, 4, 43, 1, 1, 43, 2, 11, 275, 0, 4, 
/* out0246_had-eta6-phi12*/	5, 31, 0, 6, 32, 1, 10, 42, 2, 10, 274, 0, 2, 275, 0, 1, 
/* out0247_had-eta7-phi12*/	5, 31, 0, 6, 31, 1, 11, 41, 2, 3, 42, 2, 1, 274, 0, 3, 
/* out0248_had-eta8-phi12*/	8, 30, 0, 11, 31, 1, 2, 41, 2, 4, 165, 0, 1, 165, 1, 11, 169, 0, 1, 225, 0, 3, 274, 0, 2, 
/* out0249_had-eta9-phi12*/	13, 30, 0, 1, 30, 1, 12, 40, 2, 2, 164, 0, 3, 164, 2, 3, 165, 0, 3, 165, 1, 5, 169, 0, 3, 169, 1, 3, 225, 0, 9, 225, 1, 4, 225, 2, 7, 274, 0, 1, 
/* out0250_had-eta10-phi12*/	10, 29, 0, 11, 40, 2, 1, 164, 1, 1, 164, 2, 12, 168, 0, 2, 169, 1, 1, 224, 0, 6, 224, 2, 1, 225, 1, 7, 225, 2, 2, 
/* out0251_had-eta11-phi12*/	11, 13, 8, 1, 29, 1, 9, 163, 0, 2, 163, 2, 4, 164, 1, 1, 164, 2, 1, 168, 0, 2, 168, 1, 3, 224, 0, 4, 224, 1, 3, 224, 2, 6, 
/* out0252_had-eta12-phi12*/	13, 7, 0, 15, 7, 1, 2, 7, 2, 2, 7, 3, 4, 13, 8, 3, 29, 1, 2, 163, 2, 9, 167, 0, 1, 168, 1, 1, 223, 0, 4, 223, 2, 1, 224, 1, 5, 224, 2, 1, 
/* out0253_had-eta13-phi12*/	12, 7, 1, 6, 7, 2, 11, 7, 6, 9, 7, 7, 4, 162, 2, 1, 163, 1, 1, 163, 2, 1, 167, 0, 3, 167, 1, 2, 223, 0, 3, 223, 1, 1, 223, 2, 5, 
/* out0254_had-eta14-phi12*/	8, 7, 4, 12, 7, 5, 4, 7, 6, 4, 7, 7, 3, 162, 2, 6, 167, 1, 2, 223, 1, 5, 223, 2, 3, 
/* out0255_had-eta15-phi12*/	10, 6, 0, 12, 6, 1, 1, 6, 2, 1, 6, 3, 4, 7, 4, 1, 162, 2, 4, 166, 0, 2, 222, 0, 4, 222, 2, 2, 223, 1, 1, 
/* out0256_had-eta16-phi12*/	8, 6, 1, 2, 6, 2, 11, 6, 6, 4, 161, 1, 1, 166, 0, 2, 166, 1, 2, 222, 0, 1, 222, 2, 4, 
/* out0257_had-eta17-phi12*/	8, 6, 4, 1, 6, 5, 2, 6, 6, 9, 6, 7, 2, 161, 1, 6, 166, 1, 2, 222, 1, 2, 222, 2, 2, 
/* out0258_had-eta18-phi12*/	5, 4, 0, 2, 6, 4, 7, 6, 5, 3, 161, 1, 1, 222, 1, 1, 
/* out0259_had-eta19-phi12*/	4, 4, 0, 5, 4, 1, 13, 4, 2, 1, 4, 3, 4, 
/* out0260_had-eta0-phi13*/	1, 277, 0, 1, 
/* out0261_had-eta1-phi13*/	1, 277, 0, 5, 
/* out0262_had-eta2-phi13*/	7, 45, 0, 10, 45, 1, 1, 58, 0, 2, 59, 0, 8, 59, 1, 16, 276, 0, 2, 277, 0, 2, 
/* out0263_had-eta3-phi13*/	8, 44, 0, 12, 44, 1, 1, 45, 1, 10, 57, 0, 1, 58, 0, 4, 58, 1, 4, 58, 2, 16, 276, 0, 4, 
/* out0264_had-eta4-phi13*/	6, 43, 0, 10, 44, 1, 13, 57, 0, 1, 57, 2, 14, 275, 0, 3, 276, 0, 2, 
/* out0265_had-eta5-phi13*/	6, 42, 0, 4, 43, 0, 4, 43, 1, 15, 43, 2, 2, 56, 2, 6, 275, 0, 4, 
/* out0266_had-eta6-phi13*/	6, 42, 0, 11, 42, 1, 10, 42, 2, 4, 56, 2, 1, 274, 0, 2, 275, 0, 1, 
/* out0267_had-eta7-phi13*/	6, 41, 0, 12, 41, 2, 3, 42, 1, 5, 42, 2, 1, 55, 2, 1, 274, 0, 3, 
/* out0268_had-eta8-phi13*/	9, 40, 0, 1, 41, 0, 1, 41, 1, 11, 41, 2, 6, 160, 2, 2, 165, 0, 7, 221, 0, 1, 221, 1, 8, 274, 0, 2, 
/* out0269_had-eta9-phi13*/	12, 40, 0, 7, 40, 2, 7, 160, 2, 6, 164, 0, 9, 165, 0, 5, 220, 0, 3, 220, 2, 2, 221, 0, 4, 221, 1, 8, 225, 0, 4, 225, 1, 3, 274, 0, 1, 
/* out0270_had-eta10-phi13*/	9, 13, 3, 1, 29, 0, 1, 40, 1, 5, 40, 2, 6, 164, 0, 4, 164, 1, 11, 220, 2, 12, 224, 0, 2, 225, 1, 2, 
/* out0271_had-eta11-phi13*/	14, 13, 2, 2, 13, 3, 10, 13, 8, 3, 13, 9, 15, 13, 10, 5, 29, 1, 1, 158, 2, 1, 163, 0, 9, 164, 1, 2, 219, 2, 2, 220, 1, 1, 220, 2, 1, 224, 0, 4, 224, 1, 5, 
/* out0272_had-eta12-phi13*/	13, 7, 0, 1, 7, 1, 1, 13, 5, 1, 13, 8, 9, 13, 9, 1, 13, 10, 9, 13, 11, 12, 163, 0, 2, 163, 1, 6, 163, 2, 2, 219, 2, 6, 223, 0, 3, 224, 1, 3, 
/* out0273_had-eta13-phi13*/	11, 7, 1, 7, 7, 7, 7, 11, 3, 2, 11, 9, 5, 13, 5, 3, 13, 11, 4, 162, 0, 5, 163, 1, 4, 219, 2, 1, 223, 0, 6, 223, 1, 3, 
/* out0274_had-eta14-phi13*/	10, 7, 4, 3, 7, 7, 2, 11, 8, 9, 11, 9, 10, 11, 10, 1, 162, 0, 4, 162, 1, 1, 162, 2, 3, 218, 2, 1, 223, 1, 6, 
/* out0275_had-eta15-phi13*/	8, 6, 0, 4, 6, 1, 2, 11, 8, 7, 11, 11, 6, 162, 1, 4, 162, 2, 2, 218, 2, 1, 222, 0, 6, 
/* out0276_had-eta16-phi13*/	8, 6, 1, 11, 6, 7, 4, 11, 11, 1, 161, 0, 3, 161, 1, 1, 162, 1, 1, 222, 0, 3, 222, 1, 3, 
/* out0277_had-eta17-phi13*/	7, 5, 8, 1, 5, 9, 1, 6, 4, 3, 6, 7, 9, 161, 0, 1, 161, 1, 7, 222, 1, 5, 
/* out0278_had-eta18-phi13*/	4, 4, 0, 1, 5, 8, 6, 6, 4, 5, 222, 1, 1, 
/* out0279_had-eta19-phi13*/	3, 4, 0, 8, 4, 1, 2, 5, 8, 2, 
/* out0280_had-eta0-phi14*/	1, 281, 0, 1, 
/* out0281_had-eta1-phi14*/	1, 281, 0, 5, 
/* out0282_had-eta2-phi14*/	7, 58, 0, 2, 59, 0, 8, 97, 0, 12, 97, 1, 5, 97, 2, 14, 280, 0, 2, 281, 0, 2, 
/* out0283_had-eta3-phi14*/	8, 57, 0, 3, 58, 0, 8, 58, 1, 12, 96, 0, 5, 96, 2, 13, 97, 1, 4, 97, 2, 2, 280, 0, 4, 
/* out0284_had-eta4-phi14*/	8, 57, 0, 11, 57, 1, 15, 57, 2, 2, 95, 2, 6, 96, 1, 1, 96, 2, 3, 279, 0, 3, 280, 0, 2, 
/* out0285_had-eta5-phi14*/	6, 56, 0, 15, 56, 1, 7, 56, 2, 7, 57, 1, 1, 95, 2, 1, 279, 0, 4, 
/* out0286_had-eta6-phi14*/	8, 42, 0, 1, 42, 1, 1, 55, 0, 10, 55, 2, 5, 56, 1, 7, 56, 2, 2, 278, 0, 2, 279, 0, 1, 
/* out0287_had-eta7-phi14*/	5, 41, 0, 3, 54, 0, 1, 55, 1, 6, 55, 2, 10, 278, 0, 3, 
/* out0288_had-eta8-phi14*/	10, 40, 0, 1, 41, 1, 5, 54, 0, 2, 54, 2, 10, 160, 0, 12, 160, 2, 1, 216, 0, 1, 216, 2, 2, 221, 0, 6, 278, 0, 2, 
/* out0289_had-eta9-phi14*/	11, 40, 0, 7, 40, 1, 3, 53, 2, 1, 54, 2, 4, 160, 0, 2, 160, 1, 10, 160, 2, 7, 216, 2, 6, 220, 0, 8, 221, 0, 5, 278, 0, 1, 
/* out0290_had-eta10-phi14*/	10, 13, 0, 5, 40, 1, 8, 53, 2, 3, 158, 0, 7, 158, 2, 7, 160, 1, 1, 164, 1, 1, 220, 0, 4, 220, 1, 11, 220, 2, 1, 
/* out0291_had-eta11-phi14*/	12, 13, 0, 11, 13, 1, 9, 13, 2, 14, 13, 3, 5, 13, 6, 1, 13, 7, 1, 158, 1, 3, 158, 2, 8, 163, 0, 2, 219, 0, 9, 219, 2, 1, 220, 1, 3, 
/* out0292_had-eta12-phi14*/	12, 13, 4, 6, 13, 5, 7, 13, 6, 15, 13, 7, 4, 13, 10, 2, 156, 0, 1, 156, 2, 4, 163, 0, 1, 163, 1, 4, 219, 0, 2, 219, 1, 4, 219, 2, 5, 
/* out0293_had-eta13-phi14*/	12, 11, 0, 6, 11, 2, 1, 11, 3, 13, 13, 4, 4, 13, 5, 5, 156, 2, 6, 162, 0, 3, 163, 1, 1, 218, 0, 3, 218, 2, 1, 219, 1, 3, 219, 2, 1, 
/* out0294_had-eta14-phi14*/	9, 11, 2, 9, 11, 3, 1, 11, 6, 2, 11, 9, 1, 11, 10, 10, 162, 0, 4, 162, 1, 3, 218, 0, 1, 218, 2, 7, 
/* out0295_had-eta15-phi14*/	7, 11, 5, 4, 11, 6, 5, 11, 10, 5, 11, 11, 6, 162, 1, 6, 218, 2, 5, 222, 0, 1, 
/* out0296_had-eta16-phi14*/	10, 5, 3, 5, 5, 9, 2, 6, 7, 1, 11, 5, 6, 11, 11, 3, 161, 0, 4, 162, 1, 1, 217, 2, 2, 222, 0, 1, 222, 1, 2, 
/* out0297_had-eta17-phi14*/	6, 5, 3, 2, 5, 9, 11, 5, 10, 1, 161, 0, 4, 217, 2, 4, 222, 1, 2, 
/* out0298_had-eta18-phi14*/	5, 5, 8, 5, 5, 9, 2, 5, 10, 3, 5, 11, 2, 217, 2, 1, 
/* out0299_had-eta19-phi14*/	3, 4, 1, 1, 5, 8, 2, 5, 11, 7, 
/* out0300_had-eta0-phi15*/	1, 281, 0, 1, 
/* out0301_had-eta1-phi15*/	1, 281, 0, 5, 
/* out0302_had-eta2-phi15*/	8, 97, 0, 4, 97, 1, 6, 110, 0, 11, 110, 1, 1, 110, 2, 8, 111, 1, 1, 280, 0, 2, 281, 0, 2, 
/* out0303_had-eta3-phi15*/	8, 96, 0, 11, 96, 1, 11, 97, 1, 1, 108, 0, 2, 108, 2, 6, 110, 1, 5, 110, 2, 8, 280, 0, 4, 
/* out0304_had-eta4-phi15*/	7, 95, 0, 16, 95, 1, 7, 95, 2, 5, 96, 1, 4, 108, 2, 6, 279, 0, 3, 280, 0, 2, 
/* out0305_had-eta5-phi15*/	7, 56, 0, 1, 56, 1, 2, 94, 0, 10, 94, 2, 6, 95, 1, 8, 95, 2, 4, 279, 0, 4, 
/* out0306_had-eta6-phi15*/	8, 55, 0, 6, 55, 1, 2, 93, 0, 2, 93, 2, 1, 94, 1, 5, 94, 2, 10, 278, 0, 2, 279, 0, 1, 
/* out0307_had-eta7-phi15*/	4, 54, 0, 4, 55, 1, 8, 93, 2, 9, 278, 0, 3, 
/* out0308_had-eta8-phi15*/	8, 54, 0, 9, 54, 1, 7, 54, 2, 2, 159, 0, 2, 160, 0, 2, 216, 0, 12, 216, 2, 1, 278, 0, 2, 
/* out0309_had-eta9-phi15*/	10, 53, 0, 7, 53, 2, 1, 54, 1, 7, 159, 0, 2, 159, 2, 10, 160, 1, 5, 216, 0, 2, 216, 1, 11, 216, 2, 7, 278, 0, 1, 
/* out0310_had-eta10-phi15*/	10, 53, 0, 3, 53, 1, 2, 53, 2, 8, 158, 0, 9, 158, 1, 3, 159, 2, 3, 214, 0, 6, 214, 2, 8, 220, 0, 1, 220, 1, 1, 
/* out0311_had-eta11-phi15*/	12, 12, 3, 4, 12, 9, 2, 13, 1, 7, 13, 7, 4, 53, 1, 2, 53, 2, 3, 156, 0, 2, 157, 2, 1, 158, 1, 10, 214, 1, 1, 214, 2, 8, 219, 0, 4, 
/* out0312_had-eta12-phi15*/	9, 12, 8, 8, 12, 9, 13, 13, 4, 5, 13, 7, 7, 156, 0, 9, 156, 2, 1, 213, 2, 3, 219, 0, 1, 219, 1, 7, 
/* out0313_had-eta13-phi15*/	10, 11, 0, 10, 11, 1, 6, 12, 8, 8, 12, 11, 3, 13, 4, 1, 156, 1, 5, 156, 2, 4, 213, 2, 2, 218, 0, 6, 219, 1, 2, 
/* out0314_had-eta14-phi15*/	11, 11, 1, 7, 11, 2, 6, 11, 6, 5, 11, 7, 5, 155, 0, 3, 155, 2, 2, 156, 1, 2, 156, 2, 1, 218, 0, 4, 218, 1, 3, 218, 2, 1, 
/* out0315_had-eta15-phi15*/	6, 11, 4, 9, 11, 5, 4, 11, 6, 4, 11, 7, 3, 155, 2, 6, 218, 1, 6, 
/* out0316_had-eta16-phi15*/	8, 5, 0, 6, 5, 3, 6, 11, 4, 3, 11, 5, 2, 155, 2, 4, 161, 0, 1, 217, 0, 4, 217, 2, 1, 
/* out0317_had-eta17-phi15*/	6, 5, 2, 9, 5, 3, 3, 5, 10, 2, 161, 0, 3, 217, 0, 1, 217, 2, 5, 
/* out0318_had-eta18-phi15*/	5, 5, 2, 1, 5, 6, 3, 5, 10, 8, 5, 11, 3, 217, 2, 3, 
/* out0319_had-eta19-phi15*/	4, 5, 5, 3, 5, 6, 2, 5, 10, 2, 5, 11, 4, 
/* out0320_had-eta0-phi16*/	1, 285, 0, 1, 
/* out0321_had-eta1-phi16*/	1, 285, 0, 5, 
/* out0322_had-eta2-phi16*/	8, 109, 0, 10, 109, 2, 3, 110, 0, 5, 110, 1, 4, 111, 0, 16, 111, 1, 15, 284, 0, 2, 285, 0, 2, 
/* out0323_had-eta3-phi16*/	9, 107, 0, 1, 107, 2, 2, 108, 0, 14, 108, 1, 5, 108, 2, 1, 109, 1, 4, 109, 2, 13, 110, 1, 6, 284, 0, 4, 
/* out0324_had-eta4-phi16*/	9, 95, 1, 1, 106, 0, 14, 106, 1, 1, 106, 2, 5, 107, 2, 4, 108, 1, 11, 108, 2, 3, 283, 0, 3, 284, 0, 2, 
/* out0325_had-eta5-phi16*/	7, 94, 0, 6, 94, 1, 3, 105, 0, 3, 105, 2, 2, 106, 1, 7, 106, 2, 11, 283, 0, 4, 
/* out0326_had-eta6-phi16*/	5, 93, 0, 9, 94, 1, 8, 105, 2, 9, 282, 0, 2, 283, 0, 1, 
/* out0327_had-eta7-phi16*/	4, 93, 0, 5, 93, 1, 11, 93, 2, 5, 282, 0, 3, 
/* out0328_had-eta8-phi16*/	11, 54, 1, 2, 92, 0, 7, 92, 2, 6, 93, 1, 2, 93, 2, 1, 159, 0, 4, 215, 0, 3, 215, 2, 1, 216, 0, 1, 216, 1, 1, 282, 0, 2, 
/* out0329_had-eta9-phi16*/	10, 53, 0, 4, 92, 2, 10, 159, 0, 8, 159, 1, 9, 159, 2, 2, 214, 0, 1, 215, 0, 3, 215, 2, 12, 216, 1, 4, 282, 0, 1, 
/* out0330_had-eta10-phi16*/	10, 53, 0, 2, 53, 1, 8, 132, 2, 1, 157, 0, 7, 157, 2, 2, 159, 1, 6, 159, 2, 1, 214, 0, 9, 214, 1, 6, 215, 2, 2, 
/* out0331_had-eta11-phi16*/	10, 12, 0, 13, 12, 1, 1, 12, 2, 1, 12, 3, 10, 53, 1, 4, 157, 0, 1, 157, 1, 1, 157, 2, 11, 213, 0, 4, 214, 1, 9, 
/* out0332_had-eta12-phi16*/	13, 12, 2, 13, 12, 3, 2, 12, 6, 6, 12, 9, 1, 12, 10, 13, 156, 0, 4, 156, 1, 3, 157, 1, 1, 157, 2, 2, 194, 2, 1, 213, 0, 6, 213, 1, 1, 213, 2, 5, 
/* out0333_had-eta13-phi16*/	9, 12, 5, 9, 12, 6, 3, 12, 10, 3, 12, 11, 12, 156, 1, 6, 194, 2, 2, 213, 1, 2, 213, 2, 6, 218, 0, 1, 
/* out0334_had-eta14-phi16*/	10, 11, 1, 3, 11, 7, 7, 12, 5, 1, 12, 11, 1, 16, 3, 3, 16, 9, 8, 155, 0, 7, 207, 2, 2, 218, 0, 1, 218, 1, 4, 
/* out0335_had-eta15-phi16*/	10, 11, 4, 4, 11, 7, 1, 16, 8, 9, 16, 9, 3, 155, 0, 2, 155, 1, 2, 155, 2, 2, 207, 2, 2, 217, 0, 1, 218, 1, 3, 
/* out0336_had-eta16-phi16*/	6, 5, 0, 10, 5, 1, 2, 16, 8, 4, 155, 1, 4, 155, 2, 2, 217, 0, 5, 
/* out0337_had-eta17-phi16*/	6, 5, 1, 6, 5, 2, 6, 5, 6, 1, 155, 1, 1, 217, 0, 2, 217, 1, 3, 
/* out0338_had-eta18-phi16*/	4, 5, 5, 7, 5, 6, 9, 5, 7, 2, 217, 1, 3, 
/* out0339_had-eta19-phi16*/	3, 5, 4, 3, 5, 5, 6, 5, 6, 1, 
/* out0340_had-eta0-phi17*/	1, 285, 0, 1, 
/* out0341_had-eta1-phi17*/	1, 285, 0, 5, 
/* out0342_had-eta2-phi17*/	6, 109, 0, 6, 109, 1, 2, 121, 0, 6, 121, 2, 2, 284, 0, 2, 285, 0, 2, 
/* out0343_had-eta3-phi17*/	7, 107, 0, 15, 107, 1, 3, 107, 2, 2, 109, 1, 10, 121, 0, 1, 121, 2, 14, 284, 0, 4, 
/* out0344_had-eta4-phi17*/	8, 106, 0, 2, 106, 1, 3, 107, 1, 13, 107, 2, 8, 117, 0, 8, 117, 2, 3, 283, 0, 3, 284, 0, 2, 
/* out0345_had-eta5-phi17*/	5, 105, 0, 12, 105, 1, 1, 106, 1, 5, 117, 2, 13, 283, 0, 4, 
/* out0346_had-eta6-phi17*/	6, 105, 0, 1, 105, 1, 15, 105, 2, 5, 127, 0, 3, 282, 0, 2, 283, 0, 1, 
/* out0347_had-eta7-phi17*/	4, 93, 1, 3, 127, 0, 4, 127, 2, 13, 282, 0, 3, 
/* out0348_had-eta8-phi17*/	6, 92, 0, 9, 92, 1, 5, 127, 2, 3, 197, 0, 1, 215, 0, 2, 282, 0, 2, 
/* out0349_had-eta9-phi17*/	9, 92, 1, 11, 132, 0, 3, 159, 1, 1, 197, 0, 7, 197, 2, 9, 215, 0, 8, 215, 1, 13, 215, 2, 1, 282, 0, 1, 
/* out0350_had-eta10-phi17*/	8, 132, 0, 4, 132, 2, 8, 157, 0, 7, 157, 1, 1, 197, 2, 7, 211, 0, 8, 211, 2, 5, 215, 1, 3, 
/* out0351_had-eta11-phi17*/	7, 12, 0, 3, 12, 1, 9, 132, 2, 7, 157, 0, 1, 157, 1, 11, 211, 2, 11, 213, 0, 2, 
/* out0352_had-eta12-phi17*/	10, 12, 1, 6, 12, 2, 2, 12, 4, 3, 12, 6, 6, 12, 7, 16, 157, 1, 2, 194, 0, 7, 194, 2, 1, 213, 0, 4, 213, 1, 6, 
/* out0353_had-eta13-phi17*/	9, 12, 4, 13, 12, 5, 6, 12, 6, 1, 16, 0, 6, 16, 3, 1, 194, 0, 1, 194, 2, 8, 207, 0, 2, 213, 1, 7, 
/* out0354_had-eta14-phi17*/	9, 16, 0, 1, 16, 2, 7, 16, 3, 12, 16, 9, 2, 16, 10, 2, 155, 0, 3, 194, 2, 4, 207, 0, 5, 207, 2, 3, 
/* out0355_had-eta15-phi17*/	7, 16, 8, 1, 16, 9, 3, 16, 10, 13, 16, 11, 2, 155, 0, 1, 155, 1, 5, 207, 2, 7, 
/* out0356_had-eta16-phi17*/	7, 5, 1, 2, 16, 8, 2, 16, 11, 13, 155, 1, 4, 207, 2, 2, 217, 0, 3, 217, 1, 1, 
/* out0357_had-eta17-phi17*/	3, 5, 1, 6, 5, 7, 7, 217, 1, 5, 
/* out0358_had-eta18-phi17*/	3, 5, 4, 4, 5, 7, 7, 217, 1, 4, 
/* out0359_had-eta19-phi17*/	1, 5, 4, 9, 
/* out0360_had-eta0-phi18*/	1, 289, 0, 1, 
/* out0361_had-eta1-phi18*/	1, 289, 0, 5, 
/* out0362_had-eta2-phi18*/	6, 119, 0, 6, 119, 2, 2, 121, 0, 7, 121, 1, 2, 288, 0, 2, 289, 0, 2, 
/* out0363_had-eta3-phi18*/	7, 118, 0, 15, 118, 1, 2, 118, 2, 3, 119, 2, 10, 121, 0, 2, 121, 1, 14, 288, 0, 4, 
/* out0364_had-eta4-phi18*/	8, 117, 0, 8, 117, 1, 3, 118, 1, 8, 118, 2, 13, 129, 0, 2, 129, 2, 3, 287, 0, 3, 288, 0, 2, 
/* out0365_had-eta5-phi18*/	5, 117, 1, 13, 128, 0, 12, 128, 2, 1, 129, 2, 5, 287, 0, 4, 
/* out0366_had-eta6-phi18*/	6, 127, 0, 4, 128, 0, 1, 128, 1, 5, 128, 2, 15, 286, 0, 2, 287, 0, 1, 
/* out0367_had-eta7-phi18*/	4, 127, 0, 5, 127, 1, 13, 134, 2, 3, 286, 0, 3, 
/* out0368_had-eta8-phi18*/	6, 127, 1, 3, 133, 0, 9, 133, 2, 5, 197, 0, 1, 212, 0, 2, 286, 0, 2, 
/* out0369_had-eta9-phi18*/	9, 132, 0, 4, 133, 2, 11, 196, 2, 1, 197, 0, 7, 197, 1, 9, 212, 0, 8, 212, 1, 1, 212, 2, 13, 286, 0, 1, 
/* out0370_had-eta10-phi18*/	8, 132, 0, 5, 132, 1, 7, 195, 0, 7, 195, 2, 1, 197, 1, 7, 211, 0, 8, 211, 1, 5, 212, 2, 3, 
/* out0371_had-eta11-phi18*/	7, 17, 0, 3, 17, 3, 9, 132, 1, 7, 195, 0, 1, 195, 2, 11, 208, 0, 2, 211, 1, 11, 
/* out0372_had-eta12-phi18*/	10, 17, 2, 2, 17, 3, 6, 17, 8, 3, 17, 9, 16, 17, 10, 6, 194, 0, 7, 194, 1, 1, 195, 2, 2, 208, 0, 4, 208, 2, 6, 
/* out0373_had-eta13-phi18*/	9, 16, 0, 7, 16, 1, 1, 17, 8, 13, 17, 10, 1, 17, 11, 6, 194, 0, 1, 194, 1, 8, 207, 0, 3, 208, 2, 7, 
/* out0374_had-eta14-phi18*/	9, 16, 0, 2, 16, 1, 11, 16, 2, 8, 16, 6, 2, 16, 7, 1, 151, 0, 3, 194, 1, 3, 207, 0, 5, 207, 1, 2, 
/* out0375_had-eta15-phi18*/	9, 16, 2, 1, 16, 4, 1, 16, 5, 2, 16, 6, 14, 16, 7, 2, 16, 10, 1, 151, 0, 1, 151, 2, 5, 207, 1, 6, 
/* out0376_had-eta16-phi18*/	7, 16, 5, 13, 16, 11, 1, 21, 3, 2, 151, 2, 4, 202, 0, 3, 202, 2, 1, 207, 1, 2, 
/* out0377_had-eta17-phi18*/	4, 16, 5, 1, 21, 3, 6, 21, 9, 7, 202, 2, 5, 
/* out0378_had-eta18-phi18*/	3, 21, 8, 4, 21, 9, 7, 202, 2, 4, 
/* out0379_had-eta19-phi18*/	1, 21, 8, 9, 
/* out0380_had-eta0-phi19*/	1, 289, 0, 1, 
/* out0381_had-eta1-phi19*/	1, 289, 0, 5, 
/* out0382_had-eta2-phi19*/	8, 119, 0, 10, 119, 1, 3, 120, 0, 15, 120, 1, 16, 131, 0, 5, 131, 2, 4, 288, 0, 2, 289, 0, 2, 
/* out0383_had-eta3-phi19*/	9, 118, 0, 1, 118, 1, 2, 119, 1, 13, 119, 2, 4, 130, 0, 14, 130, 1, 1, 130, 2, 5, 131, 2, 6, 288, 0, 4, 
/* out0384_had-eta4-phi19*/	9, 118, 1, 4, 129, 0, 14, 129, 1, 5, 129, 2, 1, 130, 1, 3, 130, 2, 11, 136, 2, 1, 287, 0, 3, 288, 0, 2, 
/* out0385_had-eta5-phi19*/	7, 128, 0, 3, 128, 1, 2, 129, 1, 11, 129, 2, 7, 135, 0, 6, 135, 2, 3, 287, 0, 4, 
/* out0386_had-eta6-phi19*/	5, 128, 1, 9, 134, 0, 9, 135, 2, 8, 286, 0, 2, 287, 0, 1, 
/* out0387_had-eta7-phi19*/	4, 134, 0, 5, 134, 1, 5, 134, 2, 11, 286, 0, 3, 
/* out0388_had-eta8-phi19*/	11, 68, 2, 2, 133, 0, 7, 133, 1, 6, 134, 1, 1, 134, 2, 2, 196, 0, 4, 210, 0, 1, 210, 2, 1, 212, 0, 3, 212, 1, 1, 286, 0, 2, 
/* out0389_had-eta9-phi19*/	10, 67, 0, 4, 133, 1, 10, 196, 0, 8, 196, 1, 2, 196, 2, 9, 209, 0, 1, 210, 2, 4, 212, 0, 3, 212, 1, 12, 286, 0, 1, 
/* out0390_had-eta10-phi19*/	10, 67, 0, 2, 67, 2, 8, 132, 1, 1, 195, 0, 7, 195, 1, 2, 196, 1, 1, 196, 2, 6, 209, 0, 9, 209, 2, 6, 212, 1, 2, 
/* out0391_had-eta11-phi19*/	11, 17, 0, 13, 17, 1, 10, 17, 2, 1, 17, 3, 1, 67, 2, 4, 132, 1, 1, 195, 0, 1, 195, 1, 11, 195, 2, 1, 208, 0, 4, 209, 2, 9, 
/* out0392_had-eta12-phi19*/	13, 17, 1, 2, 17, 2, 13, 17, 6, 13, 17, 7, 1, 17, 10, 6, 152, 0, 4, 152, 2, 3, 194, 1, 1, 195, 1, 2, 195, 2, 1, 208, 0, 6, 208, 1, 5, 208, 2, 1, 
/* out0393_had-eta13-phi19*/	9, 17, 5, 12, 17, 6, 3, 17, 10, 3, 17, 11, 9, 152, 2, 6, 194, 1, 3, 203, 0, 1, 208, 1, 6, 208, 2, 2, 
/* out0394_had-eta14-phi19*/	11, 16, 1, 4, 16, 7, 9, 17, 5, 1, 17, 11, 1, 22, 3, 3, 22, 9, 7, 151, 0, 7, 203, 0, 1, 203, 2, 4, 207, 0, 1, 207, 1, 3, 
/* out0395_had-eta15-phi19*/	10, 16, 4, 10, 16, 7, 4, 22, 8, 4, 22, 9, 1, 151, 0, 2, 151, 1, 2, 151, 2, 2, 202, 0, 1, 203, 2, 3, 207, 1, 3, 
/* out0396_had-eta16-phi19*/	6, 16, 4, 5, 21, 0, 10, 21, 3, 2, 151, 1, 2, 151, 2, 4, 202, 0, 5, 
/* out0397_had-eta17-phi19*/	6, 21, 2, 6, 21, 3, 6, 21, 10, 1, 151, 2, 1, 202, 0, 2, 202, 2, 3, 
/* out0398_had-eta18-phi19*/	4, 21, 9, 2, 21, 10, 9, 21, 11, 7, 202, 2, 3, 
/* out0399_had-eta19-phi19*/	3, 21, 8, 3, 21, 10, 1, 21, 11, 6, 
/* out0400_had-eta0-phi20*/	1, 293, 0, 1, 
/* out0401_had-eta1-phi20*/	1, 293, 0, 5, 
/* out0402_had-eta2-phi20*/	8, 120, 0, 1, 131, 0, 11, 131, 1, 8, 131, 2, 1, 138, 0, 4, 138, 2, 6, 292, 0, 2, 293, 0, 2, 
/* out0403_had-eta3-phi20*/	8, 130, 0, 2, 130, 1, 6, 131, 1, 8, 131, 2, 5, 137, 0, 11, 137, 2, 11, 138, 2, 1, 292, 0, 4, 
/* out0404_had-eta4-phi20*/	7, 130, 1, 6, 136, 0, 16, 136, 1, 5, 136, 2, 7, 137, 2, 4, 291, 0, 3, 292, 0, 2, 
/* out0405_had-eta5-phi20*/	7, 70, 0, 1, 70, 2, 2, 135, 0, 10, 135, 1, 6, 136, 1, 4, 136, 2, 8, 291, 0, 4, 
/* out0406_had-eta6-phi20*/	8, 69, 0, 6, 69, 2, 2, 134, 0, 2, 134, 1, 1, 135, 1, 10, 135, 2, 5, 290, 0, 2, 291, 0, 1, 
/* out0407_had-eta7-phi20*/	4, 68, 0, 4, 69, 2, 8, 134, 1, 9, 290, 0, 3, 
/* out0408_had-eta8-phi20*/	8, 68, 0, 9, 68, 1, 2, 68, 2, 7, 154, 0, 2, 196, 0, 2, 210, 0, 12, 210, 1, 1, 290, 0, 2, 
/* out0409_had-eta9-phi20*/	10, 67, 0, 7, 67, 1, 1, 68, 2, 7, 154, 2, 5, 196, 0, 2, 196, 1, 10, 210, 0, 2, 210, 1, 7, 210, 2, 11, 290, 0, 1, 
/* out0410_had-eta10-phi20*/	10, 67, 0, 3, 67, 1, 8, 67, 2, 2, 153, 0, 9, 153, 2, 3, 196, 1, 3, 205, 0, 1, 205, 2, 1, 209, 0, 6, 209, 1, 8, 
/* out0411_had-eta11-phi20*/	12, 17, 1, 4, 17, 7, 2, 23, 3, 7, 23, 9, 4, 67, 1, 3, 67, 2, 2, 152, 0, 2, 153, 2, 10, 195, 1, 1, 204, 0, 4, 209, 1, 8, 209, 2, 1, 
/* out0412_had-eta12-phi20*/	9, 17, 4, 8, 17, 7, 13, 23, 8, 5, 23, 9, 7, 152, 0, 9, 152, 1, 1, 204, 0, 1, 204, 2, 7, 208, 1, 3, 
/* out0413_had-eta13-phi20*/	10, 17, 4, 8, 17, 5, 3, 22, 0, 10, 22, 3, 6, 23, 8, 1, 152, 1, 4, 152, 2, 5, 203, 0, 6, 204, 2, 2, 208, 1, 2, 
/* out0414_had-eta14-phi20*/	11, 22, 2, 6, 22, 3, 7, 22, 9, 5, 22, 10, 5, 151, 0, 3, 151, 1, 2, 152, 1, 1, 152, 2, 2, 203, 0, 4, 203, 1, 1, 203, 2, 3, 
/* out0415_had-eta15-phi20*/	6, 22, 8, 9, 22, 9, 3, 22, 10, 4, 22, 11, 4, 151, 1, 6, 203, 2, 6, 
/* out0416_had-eta16-phi20*/	8, 21, 0, 6, 21, 1, 6, 22, 8, 3, 22, 11, 2, 146, 0, 1, 151, 1, 4, 202, 0, 4, 202, 1, 1, 
/* out0417_had-eta17-phi20*/	6, 21, 1, 3, 21, 2, 9, 21, 6, 2, 146, 0, 3, 202, 0, 1, 202, 1, 5, 
/* out0418_had-eta18-phi20*/	5, 21, 2, 1, 21, 5, 3, 21, 6, 8, 21, 10, 3, 202, 1, 3, 
/* out0419_had-eta19-phi20*/	4, 21, 5, 4, 21, 6, 2, 21, 10, 2, 21, 11, 3, 
/* out0420_had-eta0-phi21*/	1, 293, 0, 1, 
/* out0421_had-eta1-phi21*/	1, 293, 0, 5, 
/* out0422_had-eta2-phi21*/	7, 72, 0, 2, 73, 1, 8, 138, 0, 12, 138, 1, 14, 138, 2, 5, 292, 0, 2, 293, 0, 2, 
/* out0423_had-eta3-phi21*/	8, 71, 0, 3, 72, 0, 8, 72, 2, 12, 137, 0, 5, 137, 1, 13, 138, 1, 2, 138, 2, 4, 292, 0, 4, 
/* out0424_had-eta4-phi21*/	8, 71, 0, 11, 71, 1, 2, 71, 2, 15, 136, 1, 6, 137, 1, 3, 137, 2, 1, 291, 0, 3, 292, 0, 2, 
/* out0425_had-eta5-phi21*/	6, 70, 0, 15, 70, 1, 7, 70, 2, 7, 71, 2, 1, 136, 1, 1, 291, 0, 4, 
/* out0426_had-eta6-phi21*/	8, 69, 0, 10, 69, 1, 5, 70, 1, 2, 70, 2, 7, 82, 0, 1, 82, 2, 1, 290, 0, 2, 291, 0, 1, 
/* out0427_had-eta7-phi21*/	5, 68, 0, 1, 69, 1, 10, 69, 2, 6, 81, 0, 3, 290, 0, 3, 
/* out0428_had-eta8-phi21*/	10, 68, 0, 2, 68, 1, 10, 80, 0, 1, 81, 2, 5, 154, 0, 12, 154, 1, 1, 206, 1, 6, 210, 0, 1, 210, 1, 2, 290, 0, 2, 
/* out0429_had-eta9-phi21*/	11, 67, 1, 1, 68, 1, 4, 80, 0, 7, 80, 2, 3, 154, 0, 2, 154, 1, 7, 154, 2, 10, 205, 0, 8, 206, 1, 5, 210, 1, 6, 290, 0, 1, 
/* out0430_had-eta10-phi21*/	10, 23, 0, 5, 67, 1, 3, 80, 2, 8, 149, 2, 1, 153, 0, 7, 153, 1, 7, 154, 2, 1, 205, 0, 4, 205, 1, 1, 205, 2, 11, 
/* out0431_had-eta11-phi21*/	12, 23, 0, 11, 23, 1, 5, 23, 2, 14, 23, 3, 9, 23, 9, 1, 23, 10, 1, 148, 0, 2, 153, 1, 8, 153, 2, 3, 204, 0, 9, 204, 1, 1, 205, 2, 3, 
/* out0432_had-eta12-phi21*/	12, 23, 6, 2, 23, 8, 6, 23, 9, 4, 23, 10, 15, 23, 11, 7, 148, 0, 1, 148, 2, 4, 152, 0, 1, 152, 1, 4, 204, 0, 2, 204, 1, 5, 204, 2, 4, 
/* out0433_had-eta13-phi21*/	12, 22, 0, 6, 22, 1, 13, 22, 2, 1, 23, 8, 4, 23, 11, 5, 147, 0, 3, 148, 2, 1, 152, 1, 6, 203, 0, 3, 203, 1, 1, 204, 1, 1, 204, 2, 3, 
/* out0434_had-eta14-phi21*/	9, 22, 1, 1, 22, 2, 9, 22, 6, 10, 22, 7, 1, 22, 10, 2, 147, 0, 4, 147, 2, 3, 203, 0, 1, 203, 1, 7, 
/* out0435_had-eta15-phi21*/	7, 22, 5, 6, 22, 6, 5, 22, 10, 5, 22, 11, 4, 147, 2, 6, 198, 0, 1, 203, 1, 5, 
/* out0436_had-eta16-phi21*/	9, 21, 1, 5, 21, 7, 2, 22, 5, 3, 22, 11, 6, 146, 0, 4, 147, 2, 1, 198, 0, 1, 198, 2, 2, 202, 1, 2, 
/* out0437_had-eta17-phi21*/	6, 21, 1, 2, 21, 6, 1, 21, 7, 11, 146, 0, 4, 198, 2, 2, 202, 1, 4, 
/* out0438_had-eta18-phi21*/	5, 21, 4, 5, 21, 5, 2, 21, 6, 3, 21, 7, 2, 202, 1, 1, 
/* out0439_had-eta19-phi21*/	2, 21, 4, 2, 21, 5, 7, 
/* out0440_had-eta0-phi22*/	1, 297, 0, 1, 
/* out0441_had-eta1-phi22*/	1, 297, 0, 5, 
/* out0442_had-eta2-phi22*/	7, 72, 0, 2, 73, 0, 16, 73, 1, 8, 85, 0, 10, 85, 2, 1, 296, 0, 2, 297, 0, 2, 
/* out0443_had-eta3-phi22*/	8, 71, 0, 1, 72, 0, 4, 72, 1, 16, 72, 2, 4, 84, 0, 12, 84, 2, 1, 85, 2, 10, 296, 0, 4, 
/* out0444_had-eta4-phi22*/	6, 71, 0, 1, 71, 1, 14, 83, 0, 10, 84, 2, 13, 295, 0, 3, 296, 0, 2, 
/* out0445_had-eta5-phi22*/	6, 70, 1, 6, 82, 0, 4, 83, 0, 4, 83, 1, 2, 83, 2, 15, 295, 0, 4, 
/* out0446_had-eta6-phi22*/	6, 70, 1, 1, 82, 0, 11, 82, 1, 4, 82, 2, 10, 294, 0, 2, 295, 0, 1, 
/* out0447_had-eta7-phi22*/	6, 69, 1, 1, 81, 0, 12, 81, 1, 3, 82, 1, 1, 82, 2, 5, 294, 0, 3, 
/* out0448_had-eta8-phi22*/	9, 80, 0, 1, 81, 0, 1, 81, 1, 6, 81, 2, 11, 150, 1, 7, 154, 1, 2, 206, 0, 8, 206, 1, 1, 294, 0, 2, 
/* out0449_had-eta9-phi22*/	12, 80, 0, 7, 80, 1, 7, 149, 0, 9, 150, 1, 5, 154, 1, 6, 201, 0, 4, 201, 2, 3, 205, 0, 3, 205, 1, 2, 206, 0, 8, 206, 1, 4, 294, 0, 1, 
/* out0450_had-eta10-phi22*/	8, 23, 1, 1, 80, 1, 6, 80, 2, 5, 149, 0, 4, 149, 2, 11, 200, 0, 2, 201, 2, 2, 205, 1, 12, 
/* out0451_had-eta11-phi22*/	13, 23, 1, 10, 23, 2, 2, 23, 4, 3, 23, 6, 5, 23, 7, 15, 148, 0, 9, 149, 2, 2, 153, 1, 1, 200, 0, 4, 200, 2, 5, 204, 1, 2, 205, 1, 1, 205, 2, 1, 
/* out0452_had-eta12-phi22*/	11, 23, 4, 9, 23, 5, 12, 23, 6, 9, 23, 7, 1, 23, 11, 1, 148, 0, 2, 148, 1, 2, 148, 2, 6, 199, 0, 3, 200, 2, 3, 204, 1, 6, 
/* out0453_had-eta13-phi22*/	9, 22, 1, 2, 22, 7, 5, 23, 5, 4, 23, 11, 3, 147, 0, 5, 148, 2, 4, 199, 0, 6, 199, 2, 3, 204, 1, 1, 
/* out0454_had-eta14-phi22*/	8, 22, 4, 9, 22, 6, 1, 22, 7, 10, 147, 0, 4, 147, 1, 3, 147, 2, 1, 199, 2, 6, 203, 1, 1, 
/* out0455_had-eta15-phi22*/	6, 22, 4, 7, 22, 5, 6, 147, 1, 2, 147, 2, 4, 198, 0, 6, 203, 1, 1, 
/* out0456_had-eta16-phi22*/	6, 22, 5, 1, 146, 0, 3, 146, 1, 1, 147, 2, 1, 198, 0, 3, 198, 2, 3, 
/* out0457_had-eta17-phi22*/	5, 21, 4, 1, 21, 7, 1, 146, 0, 1, 146, 1, 7, 198, 2, 5, 
/* out0458_had-eta18-phi22*/	2, 21, 4, 6, 198, 2, 1, 
/* out0459_had-eta19-phi22*/	1, 21, 4, 2, 
/* out0460_had-eta0-phi23*/	1, 297, 0, 1, 
/* out0461_had-eta1-phi23*/	1, 297, 0, 5, 
/* out0462_had-eta2-phi23*/	4, 85, 0, 6, 85, 1, 8, 296, 0, 2, 297, 0, 2, 
/* out0463_had-eta3-phi23*/	5, 84, 0, 4, 84, 1, 7, 85, 1, 8, 85, 2, 5, 296, 0, 4, 
/* out0464_had-eta4-phi23*/	6, 83, 0, 2, 83, 1, 3, 84, 1, 9, 84, 2, 2, 295, 0, 3, 296, 0, 2, 
/* out0465_had-eta5-phi23*/	3, 83, 1, 11, 83, 2, 1, 295, 0, 4, 
/* out0466_had-eta6-phi23*/	3, 82, 1, 10, 294, 0, 2, 295, 0, 1, 
/* out0467_had-eta7-phi23*/	3, 81, 1, 3, 82, 1, 1, 294, 0, 3, 
/* out0468_had-eta8-phi23*/	6, 81, 1, 4, 150, 0, 11, 150, 1, 1, 201, 0, 3, 201, 1, 7, 294, 0, 2, 
/* out0469_had-eta9-phi23*/	9, 80, 1, 2, 149, 0, 3, 149, 1, 3, 150, 0, 5, 150, 1, 3, 201, 0, 9, 201, 1, 7, 201, 2, 4, 294, 0, 1, 
/* out0470_had-eta10-phi23*/	7, 80, 1, 1, 149, 1, 12, 149, 2, 1, 200, 0, 6, 200, 1, 7, 201, 1, 2, 201, 2, 7, 
/* out0471_had-eta11-phi23*/	8, 23, 4, 1, 148, 0, 2, 148, 1, 4, 149, 1, 1, 149, 2, 1, 200, 0, 4, 200, 1, 7, 200, 2, 3, 
/* out0472_had-eta12-phi23*/	6, 23, 4, 3, 148, 1, 9, 199, 0, 4, 199, 1, 1, 200, 1, 2, 200, 2, 5, 
/* out0473_had-eta13-phi23*/	6, 147, 1, 1, 148, 1, 1, 148, 2, 1, 199, 0, 3, 199, 1, 6, 199, 2, 1, 
/* out0474_had-eta14-phi23*/	3, 147, 1, 6, 199, 1, 3, 199, 2, 5, 
/* out0475_had-eta15-phi23*/	5, 147, 1, 4, 198, 0, 4, 198, 1, 2, 199, 1, 6, 199, 2, 1, 
/* out0476_had-eta16-phi23*/	3, 146, 1, 1, 198, 0, 1, 198, 1, 5, 
/* out0477_had-eta17-phi23*/	3, 146, 1, 6, 198, 1, 3, 198, 2, 2, 
/* out0478_had-eta18-phi23*/	3, 146, 1, 1, 198, 1, 6, 198, 2, 1, 
/* out0479_had-eta19-phi23*/	0, 
};