parameter integer matrixH [0:4497] = {
/* num inputs = 133(in0-in132) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1339 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	1, 110, 0, 2, 
/* out0002_had-eta2-phi0*/	1, 110, 0, 6, 
/* out0003_had-eta3-phi0*/	1, 109, 0, 5, 
/* out0004_had-eta4-phi0*/	1, 109, 0, 3, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	3, 58, 1, 1, 63, 0, 1, 63, 2, 8, 
/* out0007_had-eta7-phi0*/	3, 63, 0, 10, 63, 1, 8, 63, 2, 8, 
/* out0008_had-eta8-phi0*/	3, 62, 0, 4, 62, 2, 12, 63, 1, 8, 
/* out0009_had-eta9-phi0*/	4, 61, 2, 2, 62, 0, 3, 62, 1, 15, 62, 2, 4, 
/* out0010_had-eta10-phi0*/	3, 61, 0, 2, 61, 1, 1, 61, 2, 11, 
/* out0011_had-eta11-phi0*/	4, 60, 2, 1, 61, 0, 1, 61, 1, 14, 104, 2, 8, 
/* out0012_had-eta12-phi0*/	4, 60, 2, 10, 104, 0, 3, 104, 1, 6, 104, 2, 5, 
/* out0013_had-eta13-phi0*/	5, 60, 0, 1, 60, 1, 7, 60, 2, 1, 103, 2, 5, 104, 1, 9, 
/* out0014_had-eta14-phi0*/	5, 59, 2, 4, 60, 1, 6, 103, 0, 1, 103, 1, 3, 103, 2, 7, 
/* out0015_had-eta15-phi0*/	3, 59, 1, 1, 59, 2, 6, 103, 1, 8, 
/* out0016_had-eta16-phi0*/	3, 59, 1, 5, 102, 2, 7, 103, 1, 1, 
/* out0017_had-eta17-phi0*/	3, 59, 1, 3, 102, 1, 3, 102, 2, 3, 
/* out0018_had-eta18-phi0*/	1, 102, 1, 5, 
/* out0019_had-eta19-phi0*/	1, 102, 1, 2, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	1, 110, 0, 2, 
/* out0022_had-eta2-phi1*/	1, 110, 0, 6, 
/* out0023_had-eta3-phi1*/	1, 109, 0, 5, 
/* out0024_had-eta4-phi1*/	1, 109, 0, 3, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	2, 58, 0, 5, 58, 1, 7, 
/* out0027_had-eta7-phi1*/	3, 57, 2, 12, 58, 1, 8, 63, 0, 5, 
/* out0028_had-eta8-phi1*/	4, 56, 2, 1, 57, 1, 13, 57, 2, 3, 62, 0, 4, 
/* out0029_had-eta9-phi1*/	5, 56, 1, 2, 56, 2, 10, 61, 2, 1, 62, 0, 5, 62, 1, 1, 
/* out0030_had-eta10-phi1*/	4, 55, 2, 1, 56, 1, 6, 61, 0, 8, 61, 2, 2, 
/* out0031_had-eta11-phi1*/	8, 55, 1, 1, 55, 2, 5, 60, 2, 3, 61, 0, 5, 61, 1, 1, 100, 1, 6, 104, 0, 2, 104, 2, 3, 
/* out0032_had-eta12-phi1*/	6, 55, 1, 2, 60, 0, 7, 60, 2, 1, 98, 2, 3, 100, 1, 2, 104, 0, 9, 
/* out0033_had-eta13-phi1*/	8, 60, 0, 7, 60, 1, 1, 98, 1, 3, 98, 2, 3, 103, 0, 2, 103, 2, 2, 104, 0, 2, 104, 1, 1, 
/* out0034_had-eta14-phi1*/	8, 54, 1, 1, 54, 2, 1, 59, 0, 2, 59, 2, 5, 60, 0, 1, 60, 1, 2, 103, 0, 9, 103, 2, 2, 
/* out0035_had-eta15-phi1*/	7, 59, 0, 5, 59, 1, 1, 59, 2, 1, 97, 2, 1, 102, 2, 2, 103, 0, 4, 103, 1, 3, 
/* out0036_had-eta16-phi1*/	5, 59, 0, 3, 59, 1, 2, 102, 0, 3, 102, 2, 3, 103, 1, 1, 
/* out0037_had-eta17-phi1*/	4, 59, 1, 3, 102, 0, 5, 102, 1, 1, 102, 2, 1, 
/* out0038_had-eta18-phi1*/	2, 102, 0, 1, 102, 1, 4, 
/* out0039_had-eta19-phi1*/	1, 102, 1, 1, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	1, 112, 0, 2, 
/* out0042_had-eta2-phi2*/	1, 112, 0, 6, 
/* out0043_had-eta3-phi2*/	1, 111, 0, 5, 
/* out0044_had-eta4-phi2*/	1, 111, 0, 3, 
/* out0045_had-eta5-phi2*/	0, 
/* out0046_had-eta6-phi2*/	2, 51, 2, 10, 58, 0, 9, 
/* out0047_had-eta7-phi2*/	6, 49, 2, 1, 51, 1, 10, 51, 2, 5, 57, 0, 8, 57, 2, 1, 58, 0, 2, 
/* out0048_had-eta8-phi2*/	6, 49, 1, 2, 49, 2, 6, 56, 0, 1, 56, 2, 1, 57, 0, 8, 57, 1, 3, 
/* out0049_had-eta9-phi2*/	4, 49, 1, 1, 56, 0, 11, 56, 1, 1, 56, 2, 4, 
/* out0050_had-eta10-phi2*/	4, 55, 0, 1, 55, 2, 4, 56, 0, 2, 56, 1, 7, 
/* out0051_had-eta11-phi2*/	5, 55, 0, 3, 55, 1, 2, 55, 2, 6, 100, 0, 13, 100, 1, 5, 
/* out0052_had-eta12-phi2*/	5, 54, 2, 1, 55, 1, 9, 98, 0, 2, 98, 2, 8, 100, 1, 3, 
/* out0053_had-eta13-phi2*/	4, 54, 2, 8, 98, 0, 2, 98, 1, 7, 98, 2, 2, 
/* out0054_had-eta14-phi2*/	4, 54, 1, 5, 54, 2, 1, 97, 2, 5, 98, 1, 4, 
/* out0055_had-eta15-phi2*/	5, 53, 2, 1, 54, 1, 2, 59, 0, 3, 97, 1, 2, 97, 2, 6, 
/* out0056_had-eta16-phi2*/	4, 53, 2, 2, 59, 0, 3, 97, 1, 5, 102, 0, 1, 
/* out0057_had-eta17-phi2*/	6, 53, 1, 1, 53, 2, 1, 59, 1, 1, 96, 2, 1, 97, 1, 1, 102, 0, 4, 
/* out0058_had-eta18-phi2*/	2, 96, 2, 3, 102, 0, 2, 
/* out0059_had-eta19-phi2*/	1, 96, 1, 1, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 112, 0, 2, 
/* out0062_had-eta2-phi3*/	1, 112, 0, 6, 
/* out0063_had-eta3-phi3*/	1, 111, 0, 5, 
/* out0064_had-eta4-phi3*/	1, 111, 0, 3, 
/* out0065_had-eta5-phi3*/	0, 
/* out0066_had-eta6-phi3*/	3, 51, 0, 6, 51, 2, 1, 52, 2, 1, 
/* out0067_had-eta7-phi3*/	6, 49, 0, 2, 49, 2, 3, 51, 0, 10, 51, 1, 6, 52, 1, 2, 52, 2, 4, 
/* out0068_had-eta8-phi3*/	3, 49, 0, 8, 49, 1, 6, 49, 2, 6, 
/* out0069_had-eta9-phi3*/	3, 48, 2, 9, 49, 1, 7, 56, 0, 2, 
/* out0070_had-eta10-phi3*/	3, 48, 1, 8, 48, 2, 5, 55, 0, 1, 
/* out0071_had-eta11-phi3*/	6, 47, 2, 2, 48, 1, 1, 55, 0, 8, 100, 0, 3, 101, 1, 1, 101, 2, 15, 
/* out0072_had-eta12-phi3*/	8, 47, 1, 1, 47, 2, 2, 54, 0, 1, 54, 2, 2, 55, 0, 3, 55, 1, 2, 98, 0, 5, 101, 1, 8, 
/* out0073_had-eta13-phi3*/	5, 54, 0, 6, 54, 2, 3, 98, 0, 7, 98, 1, 1, 99, 2, 3, 
/* out0074_had-eta14-phi3*/	7, 54, 0, 2, 54, 1, 5, 97, 0, 3, 97, 2, 3, 98, 1, 1, 99, 1, 1, 99, 2, 1, 
/* out0075_had-eta15-phi3*/	5, 53, 2, 3, 54, 1, 3, 97, 0, 5, 97, 1, 1, 97, 2, 1, 
/* out0076_had-eta16-phi3*/	2, 53, 2, 5, 97, 1, 6, 
/* out0077_had-eta17-phi3*/	3, 53, 1, 6, 53, 2, 1, 96, 2, 5, 
/* out0078_had-eta18-phi3*/	2, 96, 1, 2, 96, 2, 3, 
/* out0079_had-eta19-phi3*/	1, 96, 1, 4, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 114, 0, 2, 
/* out0082_had-eta2-phi4*/	1, 114, 0, 6, 
/* out0083_had-eta3-phi4*/	1, 113, 0, 5, 
/* out0084_had-eta4-phi4*/	1, 113, 0, 3, 
/* out0085_had-eta5-phi4*/	0, 
/* out0086_had-eta6-phi4*/	2, 52, 0, 4, 52, 2, 5, 
/* out0087_had-eta7-phi4*/	3, 52, 0, 7, 52, 1, 12, 52, 2, 6, 
/* out0088_had-eta8-phi4*/	4, 49, 0, 6, 50, 1, 1, 50, 2, 12, 52, 1, 2, 
/* out0089_had-eta9-phi4*/	4, 48, 0, 8, 48, 2, 2, 50, 1, 6, 50, 2, 1, 
/* out0090_had-eta10-phi4*/	2, 48, 0, 8, 48, 1, 6, 
/* out0091_had-eta11-phi4*/	6, 47, 0, 1, 47, 2, 9, 48, 1, 1, 101, 0, 13, 101, 1, 1, 101, 2, 1, 
/* out0092_had-eta12-phi4*/	6, 47, 1, 7, 47, 2, 3, 99, 0, 1, 99, 2, 4, 101, 0, 3, 101, 1, 6, 
/* out0093_had-eta13-phi4*/	6, 42, 2, 1, 47, 1, 3, 54, 0, 4, 99, 0, 1, 99, 1, 2, 99, 2, 8, 
/* out0094_had-eta14-phi4*/	4, 42, 2, 3, 54, 0, 3, 97, 0, 1, 99, 1, 8, 
/* out0095_had-eta15-phi4*/	5, 42, 1, 1, 53, 0, 2, 53, 2, 2, 92, 2, 2, 97, 0, 5, 
/* out0096_had-eta16-phi4*/	7, 53, 0, 4, 53, 2, 1, 92, 1, 1, 92, 2, 2, 96, 2, 1, 97, 0, 2, 97, 1, 1, 
/* out0097_had-eta17-phi4*/	4, 53, 0, 1, 53, 1, 7, 96, 0, 4, 96, 2, 2, 
/* out0098_had-eta18-phi4*/	3, 96, 0, 3, 96, 1, 2, 96, 2, 1, 
/* out0099_had-eta19-phi4*/	1, 96, 1, 5, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 114, 0, 2, 
/* out0102_had-eta2-phi5*/	1, 114, 0, 6, 
/* out0103_had-eta3-phi5*/	1, 113, 0, 5, 
/* out0104_had-eta4-phi5*/	1, 113, 0, 3, 
/* out0105_had-eta5-phi5*/	0, 
/* out0106_had-eta6-phi5*/	1, 66, 2, 3, 
/* out0107_had-eta7-phi5*/	3, 52, 0, 5, 66, 1, 5, 66, 2, 13, 
/* out0108_had-eta8-phi5*/	4, 50, 0, 14, 50, 1, 1, 50, 2, 3, 66, 1, 2, 
/* out0109_had-eta9-phi5*/	3, 50, 0, 2, 50, 1, 8, 64, 2, 7, 
/* out0110_had-eta10-phi5*/	2, 64, 1, 5, 64, 2, 9, 
/* out0111_had-eta11-phi5*/	3, 47, 0, 9, 64, 1, 3, 94, 2, 12, 
/* out0112_had-eta12-phi5*/	5, 47, 0, 6, 47, 1, 4, 94, 1, 8, 94, 2, 4, 99, 0, 2, 
/* out0113_had-eta13-phi5*/	3, 42, 2, 7, 47, 1, 1, 99, 0, 10, 
/* out0114_had-eta14-phi5*/	5, 42, 1, 2, 42, 2, 5, 92, 2, 2, 99, 0, 2, 99, 1, 5, 
/* out0115_had-eta15-phi5*/	3, 42, 1, 4, 53, 0, 1, 92, 2, 8, 
/* out0116_had-eta16-phi5*/	3, 53, 0, 5, 92, 1, 5, 92, 2, 2, 
/* out0117_had-eta17-phi5*/	4, 53, 0, 3, 53, 1, 1, 92, 1, 2, 96, 0, 3, 
/* out0118_had-eta18-phi5*/	2, 53, 1, 1, 96, 0, 4, 
/* out0119_had-eta19-phi5*/	2, 96, 0, 2, 96, 1, 2, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 116, 0, 2, 
/* out0122_had-eta2-phi6*/	1, 116, 0, 6, 
/* out0123_had-eta3-phi6*/	1, 115, 0, 5, 
/* out0124_had-eta4-phi6*/	1, 115, 0, 3, 
/* out0125_had-eta5-phi6*/	0, 
/* out0126_had-eta6-phi6*/	1, 66, 0, 3, 
/* out0127_had-eta7-phi6*/	3, 66, 0, 13, 66, 1, 6, 67, 2, 5, 
/* out0128_had-eta8-phi6*/	4, 65, 0, 3, 65, 1, 1, 65, 2, 14, 66, 1, 3, 
/* out0129_had-eta9-phi6*/	3, 64, 0, 7, 65, 1, 8, 65, 2, 2, 
/* out0130_had-eta10-phi6*/	2, 64, 0, 9, 64, 1, 5, 
/* out0131_had-eta11-phi6*/	3, 43, 2, 9, 64, 1, 3, 94, 0, 12, 
/* out0132_had-eta12-phi6*/	5, 43, 1, 4, 43, 2, 6, 93, 2, 2, 94, 0, 4, 94, 1, 8, 
/* out0133_had-eta13-phi6*/	3, 42, 0, 7, 43, 1, 1, 93, 2, 10, 
/* out0134_had-eta14-phi6*/	5, 42, 0, 4, 42, 1, 3, 92, 0, 3, 93, 1, 5, 93, 2, 2, 
/* out0135_had-eta15-phi6*/	3, 36, 2, 1, 42, 1, 5, 92, 0, 7, 
/* out0136_had-eta16-phi6*/	3, 36, 2, 5, 92, 0, 1, 92, 1, 5, 
/* out0137_had-eta17-phi6*/	4, 36, 1, 1, 36, 2, 3, 92, 1, 2, 105, 2, 3, 
/* out0138_had-eta18-phi6*/	2, 36, 1, 1, 105, 2, 4, 
/* out0139_had-eta19-phi6*/	2, 105, 1, 2, 105, 2, 2, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 116, 0, 2, 
/* out0142_had-eta2-phi7*/	1, 116, 0, 6, 
/* out0143_had-eta3-phi7*/	1, 115, 0, 5, 
/* out0144_had-eta4-phi7*/	1, 115, 0, 3, 
/* out0145_had-eta5-phi7*/	0, 
/* out0146_had-eta6-phi7*/	2, 67, 0, 5, 67, 2, 4, 
/* out0147_had-eta7-phi7*/	3, 67, 0, 6, 67, 1, 12, 67, 2, 7, 
/* out0148_had-eta8-phi7*/	4, 45, 2, 6, 65, 0, 12, 65, 1, 1, 67, 1, 2, 
/* out0149_had-eta9-phi7*/	4, 44, 0, 2, 44, 2, 8, 65, 0, 1, 65, 1, 6, 
/* out0150_had-eta10-phi7*/	2, 44, 1, 6, 44, 2, 8, 
/* out0151_had-eta11-phi7*/	6, 43, 0, 9, 43, 2, 1, 44, 1, 1, 95, 0, 1, 95, 1, 1, 95, 2, 13, 
/* out0152_had-eta12-phi7*/	6, 43, 0, 3, 43, 1, 7, 93, 0, 4, 93, 2, 1, 95, 1, 6, 95, 2, 3, 
/* out0153_had-eta13-phi7*/	6, 37, 2, 4, 42, 0, 2, 43, 1, 3, 93, 0, 8, 93, 1, 2, 93, 2, 1, 
/* out0154_had-eta14-phi7*/	4, 37, 2, 3, 42, 0, 3, 93, 1, 8, 106, 2, 1, 
/* out0155_had-eta15-phi7*/	5, 36, 0, 2, 36, 2, 2, 42, 1, 1, 92, 0, 3, 106, 2, 5, 
/* out0156_had-eta16-phi7*/	7, 36, 0, 1, 36, 2, 4, 92, 0, 2, 92, 1, 1, 105, 0, 1, 106, 1, 1, 106, 2, 2, 
/* out0157_had-eta17-phi7*/	4, 36, 1, 7, 36, 2, 1, 105, 0, 2, 105, 2, 4, 
/* out0158_had-eta18-phi7*/	3, 105, 0, 1, 105, 1, 2, 105, 2, 3, 
/* out0159_had-eta19-phi7*/	1, 105, 1, 5, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 118, 0, 2, 
/* out0162_had-eta2-phi8*/	1, 118, 0, 6, 
/* out0163_had-eta3-phi8*/	1, 117, 0, 5, 
/* out0164_had-eta4-phi8*/	1, 117, 0, 3, 
/* out0165_had-eta5-phi8*/	0, 
/* out0166_had-eta6-phi8*/	3, 46, 0, 1, 46, 2, 6, 67, 0, 1, 
/* out0167_had-eta7-phi8*/	6, 45, 0, 3, 45, 2, 2, 46, 1, 6, 46, 2, 10, 67, 0, 4, 67, 1, 2, 
/* out0168_had-eta8-phi8*/	3, 45, 0, 6, 45, 1, 6, 45, 2, 8, 
/* out0169_had-eta9-phi8*/	3, 39, 2, 2, 44, 0, 9, 45, 1, 7, 
/* out0170_had-eta10-phi8*/	3, 38, 2, 1, 44, 0, 5, 44, 1, 8, 
/* out0171_had-eta11-phi8*/	6, 38, 2, 8, 43, 0, 2, 44, 1, 1, 95, 0, 15, 95, 1, 1, 108, 1, 3, 
/* out0172_had-eta12-phi8*/	8, 37, 0, 2, 37, 2, 1, 38, 1, 2, 38, 2, 3, 43, 0, 2, 43, 1, 1, 95, 1, 8, 107, 2, 5, 
/* out0173_had-eta13-phi8*/	5, 37, 0, 3, 37, 2, 6, 93, 0, 3, 107, 1, 1, 107, 2, 7, 
/* out0174_had-eta14-phi8*/	7, 37, 1, 5, 37, 2, 2, 93, 0, 1, 93, 1, 1, 106, 0, 3, 106, 2, 3, 107, 1, 1, 
/* out0175_had-eta15-phi8*/	5, 36, 0, 3, 37, 1, 3, 106, 0, 1, 106, 1, 1, 106, 2, 5, 
/* out0176_had-eta16-phi8*/	2, 36, 0, 5, 106, 1, 6, 
/* out0177_had-eta17-phi8*/	3, 36, 0, 1, 36, 1, 6, 105, 0, 5, 
/* out0178_had-eta18-phi8*/	2, 105, 0, 3, 105, 1, 2, 
/* out0179_had-eta19-phi8*/	1, 105, 1, 4, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 118, 0, 2, 
/* out0182_had-eta2-phi9*/	1, 118, 0, 6, 
/* out0183_had-eta3-phi9*/	1, 117, 0, 5, 
/* out0184_had-eta4-phi9*/	1, 117, 0, 3, 
/* out0185_had-eta5-phi9*/	0, 
/* out0186_had-eta6-phi9*/	2, 41, 1, 9, 46, 0, 10, 
/* out0187_had-eta7-phi9*/	6, 40, 0, 1, 40, 2, 8, 41, 1, 2, 45, 0, 1, 46, 0, 5, 46, 1, 10, 
/* out0188_had-eta8-phi9*/	6, 39, 0, 1, 39, 2, 1, 40, 1, 3, 40, 2, 8, 45, 0, 6, 45, 1, 2, 
/* out0189_had-eta9-phi9*/	4, 39, 0, 4, 39, 1, 1, 39, 2, 11, 45, 1, 1, 
/* out0190_had-eta10-phi9*/	4, 38, 0, 4, 38, 2, 1, 39, 1, 7, 39, 2, 2, 
/* out0191_had-eta11-phi9*/	5, 38, 0, 6, 38, 1, 2, 38, 2, 3, 108, 0, 5, 108, 1, 13, 
/* out0192_had-eta12-phi9*/	5, 37, 0, 1, 38, 1, 9, 107, 0, 8, 107, 2, 2, 108, 0, 3, 
/* out0193_had-eta13-phi9*/	4, 37, 0, 8, 107, 0, 2, 107, 1, 7, 107, 2, 2, 
/* out0194_had-eta14-phi9*/	4, 37, 0, 1, 37, 1, 5, 106, 0, 5, 107, 1, 4, 
/* out0195_had-eta15-phi9*/	5, 31, 2, 3, 36, 0, 1, 37, 1, 2, 106, 0, 6, 106, 1, 2, 
/* out0196_had-eta16-phi9*/	4, 31, 2, 3, 36, 0, 2, 89, 2, 1, 106, 1, 5, 
/* out0197_had-eta17-phi9*/	5, 36, 0, 1, 36, 1, 1, 89, 2, 4, 105, 0, 1, 106, 1, 1, 
/* out0198_had-eta18-phi9*/	2, 89, 2, 2, 105, 0, 3, 
/* out0199_had-eta19-phi9*/	1, 105, 1, 1, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 120, 0, 2, 
/* out0202_had-eta2-phi10*/	1, 120, 0, 6, 
/* out0203_had-eta3-phi10*/	1, 119, 0, 5, 
/* out0204_had-eta4-phi10*/	1, 119, 0, 3, 
/* out0205_had-eta5-phi10*/	0, 
/* out0206_had-eta6-phi10*/	2, 41, 0, 7, 41, 1, 5, 
/* out0207_had-eta7-phi10*/	3, 35, 2, 5, 40, 0, 12, 41, 0, 8, 
/* out0208_had-eta8-phi10*/	4, 34, 2, 4, 39, 0, 1, 40, 0, 3, 40, 1, 13, 
/* out0209_had-eta9-phi10*/	3, 34, 2, 5, 39, 0, 10, 39, 1, 2, 
/* out0210_had-eta10-phi10*/	3, 33, 2, 8, 38, 0, 1, 39, 1, 6, 
/* out0211_had-eta11-phi10*/	6, 33, 1, 1, 33, 2, 5, 38, 0, 5, 38, 1, 1, 91, 2, 2, 108, 0, 6, 
/* out0212_had-eta12-phi10*/	6, 32, 0, 1, 32, 2, 7, 38, 1, 2, 91, 2, 9, 107, 0, 3, 108, 0, 2, 
/* out0213_had-eta13-phi10*/	8, 32, 1, 1, 32, 2, 7, 90, 0, 1, 90, 2, 2, 91, 1, 1, 91, 2, 2, 107, 0, 3, 107, 1, 3, 
/* out0214_had-eta14-phi10*/	7, 31, 0, 2, 31, 2, 2, 32, 1, 2, 32, 2, 1, 37, 0, 1, 37, 1, 1, 90, 2, 9, 
/* out0215_had-eta15-phi10*/	5, 31, 0, 1, 31, 2, 5, 90, 1, 2, 90, 2, 4, 106, 0, 1, 
/* out0216_had-eta16-phi10*/	4, 31, 1, 2, 31, 2, 3, 89, 0, 3, 89, 2, 3, 
/* out0217_had-eta17-phi10*/	2, 31, 1, 2, 89, 2, 5, 
/* out0218_had-eta18-phi10*/	2, 89, 1, 3, 89, 2, 1, 
/* out0219_had-eta19-phi10*/	1, 89, 1, 1, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 120, 0, 2, 
/* out0222_had-eta2-phi11*/	1, 120, 0, 6, 
/* out0223_had-eta3-phi11*/	1, 119, 0, 5, 
/* out0224_had-eta4-phi11*/	1, 119, 0, 3, 
/* out0225_had-eta5-phi11*/	0, 
/* out0226_had-eta6-phi11*/	3, 35, 0, 5, 35, 2, 1, 41, 0, 1, 
/* out0227_had-eta7-phi11*/	3, 35, 0, 7, 35, 1, 8, 35, 2, 10, 
/* out0228_had-eta8-phi11*/	3, 34, 0, 12, 34, 2, 4, 35, 1, 4, 
/* out0229_had-eta9-phi11*/	4, 33, 0, 1, 34, 0, 1, 34, 1, 12, 34, 2, 3, 
/* out0230_had-eta10-phi11*/	3, 33, 0, 11, 33, 1, 1, 33, 2, 2, 
/* out0231_had-eta11-phi11*/	3, 33, 1, 10, 33, 2, 1, 91, 0, 7, 
/* out0232_had-eta12-phi11*/	4, 32, 0, 10, 91, 0, 5, 91, 1, 5, 91, 2, 3, 
/* out0233_had-eta13-phi11*/	5, 32, 0, 1, 32, 1, 7, 32, 2, 1, 90, 0, 5, 91, 1, 6, 
/* out0234_had-eta14-phi11*/	5, 31, 0, 4, 32, 1, 3, 90, 0, 6, 90, 1, 2, 90, 2, 1, 
/* out0235_had-eta15-phi11*/	2, 31, 0, 6, 90, 1, 8, 
/* out0236_had-eta16-phi11*/	2, 31, 1, 5, 89, 0, 6, 
/* out0237_had-eta17-phi11*/	3, 31, 1, 3, 89, 0, 3, 89, 1, 2, 
/* out0238_had-eta18-phi11*/	1, 89, 1, 5, 
/* out0239_had-eta19-phi11*/	1, 89, 1, 1, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 122, 0, 2, 
/* out0242_had-eta2-phi12*/	1, 122, 0, 6, 
/* out0243_had-eta3-phi12*/	1, 121, 0, 5, 
/* out0244_had-eta4-phi12*/	1, 121, 0, 3, 
/* out0245_had-eta5-phi12*/	0, 
/* out0246_had-eta6-phi12*/	2, 30, 0, 2, 30, 1, 9, 
/* out0247_had-eta7-phi12*/	6, 29, 0, 5, 29, 2, 4, 30, 0, 5, 30, 1, 7, 35, 0, 4, 35, 1, 4, 
/* out0248_had-eta8-phi12*/	3, 29, 1, 4, 29, 2, 12, 34, 0, 3, 
/* out0249_had-eta9-phi12*/	3, 28, 0, 3, 28, 2, 9, 34, 1, 4, 
/* out0250_had-eta10-phi12*/	5, 27, 0, 1, 28, 1, 2, 28, 2, 7, 33, 0, 4, 33, 1, 1, 
/* out0251_had-eta11-phi12*/	5, 27, 0, 1, 27, 2, 8, 33, 1, 3, 88, 1, 12, 91, 0, 1, 
/* out0252_had-eta12-phi12*/	8, 27, 2, 6, 32, 0, 3, 87, 0, 1, 87, 2, 2, 88, 0, 2, 88, 1, 3, 91, 0, 3, 91, 1, 3, 
/* out0253_had-eta13-phi12*/	7, 26, 0, 1, 26, 2, 3, 32, 0, 1, 32, 1, 3, 87, 2, 9, 90, 0, 1, 91, 1, 1, 
/* out0254_had-eta14-phi12*/	5, 26, 2, 6, 87, 1, 1, 87, 2, 3, 90, 0, 3, 90, 1, 2, 
/* out0255_had-eta15-phi12*/	4, 26, 2, 2, 31, 0, 3, 86, 2, 5, 90, 1, 2, 
/* out0256_had-eta16-phi12*/	4, 25, 1, 3, 31, 1, 3, 86, 2, 5, 89, 0, 2, 
/* out0257_had-eta17-phi12*/	6, 25, 1, 4, 31, 1, 1, 85, 1, 1, 86, 2, 1, 89, 0, 2, 89, 1, 2, 
/* out0258_had-eta18-phi12*/	2, 85, 1, 5, 89, 1, 2, 
/* out0259_had-eta19-phi12*/	1, 85, 1, 2, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 122, 0, 2, 
/* out0262_had-eta2-phi13*/	1, 122, 0, 6, 
/* out0263_had-eta3-phi13*/	1, 121, 0, 5, 
/* out0264_had-eta4-phi13*/	1, 121, 0, 3, 
/* out0265_had-eta5-phi13*/	0, 
/* out0266_had-eta6-phi13*/	3, 24, 0, 2, 24, 2, 2, 30, 0, 5, 
/* out0267_had-eta7-phi13*/	3, 24, 2, 12, 29, 0, 8, 30, 0, 4, 
/* out0268_had-eta8-phi13*/	3, 23, 2, 5, 29, 0, 3, 29, 1, 12, 
/* out0269_had-eta9-phi13*/	3, 23, 2, 2, 28, 0, 12, 28, 1, 2, 
/* out0270_had-eta10-phi13*/	3, 22, 2, 1, 27, 0, 2, 28, 1, 11, 
/* out0271_had-eta11-phi13*/	5, 27, 0, 9, 27, 1, 1, 27, 2, 1, 88, 0, 9, 88, 1, 1, 
/* out0272_had-eta12-phi13*/	5, 27, 1, 9, 27, 2, 1, 84, 2, 1, 87, 0, 8, 88, 0, 4, 
/* out0273_had-eta13-phi13*/	6, 26, 0, 7, 26, 2, 1, 27, 1, 1, 87, 0, 4, 87, 1, 5, 87, 2, 2, 
/* out0274_had-eta14-phi13*/	5, 26, 0, 1, 26, 1, 2, 26, 2, 3, 86, 0, 3, 87, 1, 6, 
/* out0275_had-eta15-phi13*/	5, 25, 0, 1, 26, 1, 4, 26, 2, 1, 86, 0, 5, 86, 2, 2, 
/* out0276_had-eta16-phi13*/	4, 25, 0, 3, 25, 1, 4, 86, 1, 4, 86, 2, 3, 
/* out0277_had-eta17-phi13*/	4, 25, 1, 5, 85, 0, 3, 85, 1, 1, 86, 1, 2, 
/* out0278_had-eta18-phi13*/	2, 85, 0, 1, 85, 1, 6, 
/* out0279_had-eta19-phi13*/	1, 85, 1, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 124, 0, 2, 
/* out0282_had-eta2-phi14*/	1, 124, 0, 6, 
/* out0283_had-eta3-phi14*/	1, 123, 0, 5, 
/* out0284_had-eta4-phi14*/	1, 123, 0, 3, 
/* out0285_had-eta5-phi14*/	0, 
/* out0286_had-eta6-phi14*/	1, 24, 0, 9, 
/* out0287_had-eta7-phi14*/	5, 18, 2, 3, 23, 0, 1, 24, 0, 5, 24, 1, 16, 24, 2, 2, 
/* out0288_had-eta8-phi14*/	3, 23, 0, 13, 23, 1, 3, 23, 2, 5, 
/* out0289_had-eta9-phi14*/	6, 22, 0, 4, 22, 2, 1, 23, 1, 8, 23, 2, 4, 28, 0, 1, 28, 1, 1, 
/* out0290_had-eta10-phi14*/	3, 22, 0, 3, 22, 1, 1, 22, 2, 11, 
/* out0291_had-eta11-phi14*/	9, 21, 0, 1, 21, 2, 1, 22, 1, 2, 22, 2, 3, 27, 0, 3, 27, 1, 2, 84, 0, 7, 84, 2, 5, 88, 0, 1, 
/* out0292_had-eta12-phi14*/	5, 21, 2, 6, 27, 1, 3, 84, 1, 2, 84, 2, 10, 87, 0, 1, 
/* out0293_had-eta13-phi14*/	7, 21, 2, 3, 26, 0, 6, 82, 0, 1, 82, 2, 3, 84, 1, 1, 87, 0, 2, 87, 1, 3, 
/* out0294_had-eta14-phi14*/	5, 26, 0, 1, 26, 1, 5, 82, 2, 6, 86, 0, 2, 87, 1, 1, 
/* out0295_had-eta15-phi14*/	6, 20, 2, 1, 25, 0, 1, 26, 1, 4, 82, 2, 1, 86, 0, 6, 86, 1, 2, 
/* out0296_had-eta16-phi14*/	2, 25, 0, 5, 86, 1, 6, 
/* out0297_had-eta17-phi14*/	3, 25, 0, 2, 85, 0, 4, 86, 1, 1, 
/* out0298_had-eta18-phi14*/	1, 85, 0, 4, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 124, 0, 2, 
/* out0302_had-eta2-phi15*/	1, 124, 0, 6, 
/* out0303_had-eta3-phi15*/	1, 123, 0, 5, 
/* out0304_had-eta4-phi15*/	1, 123, 0, 3, 
/* out0305_had-eta5-phi15*/	0, 
/* out0306_had-eta6-phi15*/	2, 18, 0, 1, 19, 1, 3, 
/* out0307_had-eta7-phi15*/	3, 18, 0, 12, 18, 1, 4, 18, 2, 9, 
/* out0308_had-eta8-phi15*/	6, 16, 0, 4, 16, 2, 3, 18, 1, 5, 18, 2, 4, 23, 0, 2, 23, 1, 3, 
/* out0309_had-eta9-phi15*/	3, 16, 2, 11, 22, 0, 4, 23, 1, 2, 
/* out0310_had-eta10-phi15*/	2, 22, 0, 5, 22, 1, 8, 
/* out0311_had-eta11-phi15*/	5, 15, 2, 1, 21, 0, 6, 22, 1, 5, 84, 0, 9, 84, 1, 1, 
/* out0312_had-eta12-phi15*/	5, 21, 0, 5, 21, 1, 2, 21, 2, 3, 83, 2, 1, 84, 1, 11, 
/* out0313_had-eta13-phi15*/	6, 20, 0, 1, 21, 1, 5, 21, 2, 3, 82, 0, 10, 82, 2, 1, 84, 1, 1, 
/* out0314_had-eta14-phi15*/	6, 20, 0, 2, 20, 2, 4, 26, 1, 1, 82, 0, 1, 82, 1, 4, 82, 2, 4, 
/* out0315_had-eta15-phi15*/	6, 20, 2, 6, 81, 0, 2, 81, 2, 1, 82, 1, 3, 82, 2, 1, 86, 1, 1, 
/* out0316_had-eta16-phi15*/	3, 20, 2, 2, 25, 0, 3, 81, 2, 6, 
/* out0317_had-eta17-phi15*/	3, 25, 0, 1, 81, 2, 5, 85, 0, 1, 
/* out0318_had-eta18-phi15*/	1, 85, 0, 3, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 126, 0, 2, 
/* out0322_had-eta2-phi16*/	1, 126, 0, 6, 
/* out0323_had-eta3-phi16*/	1, 125, 0, 5, 
/* out0324_had-eta4-phi16*/	1, 125, 0, 3, 
/* out0325_had-eta5-phi16*/	0, 
/* out0326_had-eta6-phi16*/	2, 19, 0, 7, 19, 1, 10, 
/* out0327_had-eta7-phi16*/	6, 17, 0, 4, 17, 2, 6, 18, 0, 3, 18, 1, 5, 19, 0, 4, 19, 1, 3, 
/* out0328_had-eta8-phi16*/	4, 16, 0, 11, 16, 1, 1, 17, 2, 7, 18, 1, 2, 
/* out0329_had-eta9-phi16*/	4, 15, 0, 1, 16, 0, 1, 16, 1, 13, 16, 2, 2, 
/* out0330_had-eta10-phi16*/	3, 15, 0, 7, 15, 2, 6, 16, 1, 1, 
/* out0331_had-eta11-phi16*/	5, 15, 1, 2, 15, 2, 9, 21, 0, 2, 83, 0, 6, 83, 2, 1, 
/* out0332_had-eta12-phi16*/	6, 11, 2, 1, 21, 0, 2, 21, 1, 5, 83, 0, 2, 83, 1, 1, 83, 2, 10, 
/* out0333_had-eta13-phi16*/	7, 11, 2, 1, 20, 0, 3, 21, 1, 4, 82, 0, 4, 82, 1, 1, 83, 1, 1, 83, 2, 4, 
/* out0334_had-eta14-phi16*/	3, 20, 0, 7, 79, 2, 2, 82, 1, 7, 
/* out0335_had-eta15-phi16*/	5, 20, 1, 3, 20, 2, 2, 79, 2, 1, 81, 0, 6, 82, 1, 1, 
/* out0336_had-eta16-phi16*/	5, 20, 1, 3, 20, 2, 1, 81, 0, 4, 81, 1, 1, 81, 2, 1, 
/* out0337_had-eta17-phi16*/	2, 81, 1, 4, 81, 2, 2, 
/* out0338_had-eta18-phi16*/	2, 81, 1, 1, 81, 2, 1, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 126, 0, 2, 
/* out0342_had-eta2-phi17*/	1, 126, 0, 6, 
/* out0343_had-eta3-phi17*/	1, 125, 0, 5, 
/* out0344_had-eta4-phi17*/	1, 125, 0, 3, 
/* out0345_had-eta5-phi17*/	0, 
/* out0346_had-eta6-phi17*/	2, 19, 0, 4, 71, 1, 9, 
/* out0347_had-eta7-phi17*/	5, 17, 0, 12, 17, 1, 6, 17, 2, 1, 19, 0, 1, 71, 1, 7, 
/* out0348_had-eta8-phi17*/	4, 17, 1, 10, 17, 2, 2, 68, 0, 6, 68, 2, 1, 
/* out0349_had-eta9-phi17*/	4, 15, 0, 1, 16, 1, 1, 68, 0, 1, 68, 2, 13, 
/* out0350_had-eta10-phi17*/	3, 15, 0, 7, 15, 1, 5, 68, 2, 2, 
/* out0351_had-eta11-phi17*/	3, 11, 0, 2, 15, 1, 9, 83, 0, 5, 
/* out0352_had-eta12-phi17*/	4, 11, 0, 6, 11, 2, 5, 83, 0, 3, 83, 1, 10, 
/* out0353_had-eta13-phi17*/	3, 11, 2, 8, 79, 0, 6, 83, 1, 4, 
/* out0354_had-eta14-phi17*/	5, 11, 2, 1, 20, 0, 3, 20, 1, 2, 79, 0, 1, 79, 2, 8, 
/* out0355_had-eta15-phi17*/	3, 20, 1, 6, 79, 2, 5, 81, 0, 3, 
/* out0356_had-eta16-phi17*/	3, 20, 1, 2, 81, 0, 1, 81, 1, 5, 
/* out0357_had-eta17-phi17*/	1, 81, 1, 5, 
/* out0358_had-eta18-phi17*/	0, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 128, 0, 2, 
/* out0362_had-eta2-phi18*/	1, 128, 0, 6, 
/* out0363_had-eta3-phi18*/	1, 127, 0, 5, 
/* out0364_had-eta4-phi18*/	1, 127, 0, 3, 
/* out0365_had-eta5-phi18*/	0, 
/* out0366_had-eta6-phi18*/	2, 70, 1, 4, 71, 0, 9, 
/* out0367_had-eta7-phi18*/	5, 69, 0, 12, 69, 1, 1, 69, 2, 6, 70, 1, 1, 71, 0, 7, 
/* out0368_had-eta8-phi18*/	4, 68, 0, 7, 68, 1, 1, 69, 1, 2, 69, 2, 10, 
/* out0369_had-eta9-phi18*/	4, 12, 0, 1, 13, 2, 1, 68, 0, 2, 68, 1, 13, 
/* out0370_had-eta10-phi18*/	3, 12, 0, 7, 12, 2, 5, 68, 1, 2, 
/* out0371_had-eta11-phi18*/	3, 11, 0, 2, 12, 2, 9, 80, 0, 5, 
/* out0372_had-eta12-phi18*/	4, 11, 0, 6, 11, 1, 4, 80, 0, 3, 80, 2, 10, 
/* out0373_had-eta13-phi18*/	3, 11, 1, 7, 79, 0, 7, 80, 2, 4, 
/* out0374_had-eta14-phi18*/	5, 6, 0, 3, 6, 2, 2, 11, 1, 1, 79, 0, 2, 79, 1, 7, 
/* out0375_had-eta15-phi18*/	3, 6, 2, 6, 76, 0, 3, 79, 1, 5, 
/* out0376_had-eta16-phi18*/	3, 6, 2, 2, 76, 0, 1, 76, 2, 5, 
/* out0377_had-eta17-phi18*/	1, 76, 2, 5, 
/* out0378_had-eta18-phi18*/	0, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 128, 0, 2, 
/* out0382_had-eta2-phi19*/	1, 128, 0, 6, 
/* out0383_had-eta3-phi19*/	1, 127, 0, 5, 
/* out0384_had-eta4-phi19*/	1, 127, 0, 3, 
/* out0385_had-eta5-phi19*/	0, 
/* out0386_had-eta6-phi19*/	2, 70, 0, 10, 70, 1, 7, 
/* out0387_had-eta7-phi19*/	6, 14, 0, 3, 14, 2, 5, 69, 0, 4, 69, 1, 6, 70, 0, 3, 70, 1, 4, 
/* out0388_had-eta8-phi19*/	4, 13, 0, 11, 13, 2, 1, 14, 2, 2, 69, 1, 7, 
/* out0389_had-eta9-phi19*/	4, 12, 0, 1, 13, 0, 1, 13, 1, 2, 13, 2, 13, 
/* out0390_had-eta10-phi19*/	3, 12, 0, 7, 12, 1, 6, 13, 2, 1, 
/* out0391_had-eta11-phi19*/	5, 7, 0, 2, 12, 1, 9, 12, 2, 2, 80, 0, 6, 80, 1, 1, 
/* out0392_had-eta12-phi19*/	6, 7, 0, 2, 7, 2, 5, 11, 1, 2, 80, 0, 2, 80, 1, 10, 80, 2, 1, 
/* out0393_had-eta13-phi19*/	8, 6, 0, 3, 7, 2, 4, 11, 1, 2, 77, 0, 4, 77, 2, 1, 79, 1, 1, 80, 1, 4, 80, 2, 1, 
/* out0394_had-eta14-phi19*/	3, 6, 0, 7, 77, 2, 7, 79, 1, 2, 
/* out0395_had-eta15-phi19*/	5, 6, 1, 2, 6, 2, 3, 76, 0, 6, 77, 2, 1, 79, 1, 1, 
/* out0396_had-eta16-phi19*/	5, 6, 1, 1, 6, 2, 3, 76, 0, 4, 76, 1, 1, 76, 2, 1, 
/* out0397_had-eta17-phi19*/	2, 76, 1, 2, 76, 2, 4, 
/* out0398_had-eta18-phi19*/	2, 76, 1, 1, 76, 2, 1, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 130, 0, 2, 
/* out0402_had-eta2-phi20*/	1, 130, 0, 6, 
/* out0403_had-eta3-phi20*/	1, 129, 0, 5, 
/* out0404_had-eta4-phi20*/	1, 129, 0, 3, 
/* out0405_had-eta5-phi20*/	0, 
/* out0406_had-eta6-phi20*/	2, 14, 0, 1, 70, 0, 3, 
/* out0407_had-eta7-phi20*/	3, 14, 0, 12, 14, 1, 9, 14, 2, 4, 
/* out0408_had-eta8-phi20*/	6, 9, 0, 2, 9, 2, 3, 13, 0, 4, 13, 1, 3, 14, 1, 4, 14, 2, 5, 
/* out0409_had-eta9-phi20*/	3, 8, 0, 4, 9, 2, 2, 13, 1, 11, 
/* out0410_had-eta10-phi20*/	2, 8, 0, 5, 8, 2, 8, 
/* out0411_had-eta11-phi20*/	5, 7, 0, 6, 8, 2, 5, 12, 1, 1, 78, 0, 9, 78, 2, 1, 
/* out0412_had-eta12-phi20*/	5, 7, 0, 5, 7, 1, 3, 7, 2, 2, 78, 2, 11, 80, 1, 1, 
/* out0413_had-eta13-phi20*/	6, 6, 0, 1, 7, 1, 3, 7, 2, 5, 77, 0, 10, 77, 1, 1, 78, 2, 1, 
/* out0414_had-eta14-phi20*/	6, 1, 2, 1, 6, 0, 2, 6, 1, 4, 77, 0, 1, 77, 1, 4, 77, 2, 4, 
/* out0415_had-eta15-phi20*/	6, 6, 1, 6, 73, 2, 1, 76, 0, 2, 76, 1, 1, 77, 1, 1, 77, 2, 3, 
/* out0416_had-eta16-phi20*/	3, 0, 0, 3, 6, 1, 2, 76, 1, 6, 
/* out0417_had-eta17-phi20*/	3, 0, 0, 1, 72, 0, 1, 76, 1, 5, 
/* out0418_had-eta18-phi20*/	1, 72, 0, 3, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 130, 0, 2, 
/* out0422_had-eta2-phi21*/	1, 130, 0, 6, 
/* out0423_had-eta3-phi21*/	1, 129, 0, 5, 
/* out0424_had-eta4-phi21*/	1, 129, 0, 3, 
/* out0425_had-eta5-phi21*/	0, 
/* out0426_had-eta6-phi21*/	1, 10, 0, 9, 
/* out0427_had-eta7-phi21*/	5, 9, 0, 1, 10, 0, 5, 10, 1, 2, 10, 2, 16, 14, 1, 3, 
/* out0428_had-eta8-phi21*/	3, 9, 0, 13, 9, 1, 5, 9, 2, 3, 
/* out0429_had-eta9-phi21*/	6, 3, 0, 1, 3, 2, 1, 8, 0, 4, 8, 1, 1, 9, 1, 4, 9, 2, 8, 
/* out0430_had-eta10-phi21*/	3, 8, 0, 3, 8, 1, 11, 8, 2, 1, 
/* out0431_had-eta11-phi21*/	9, 2, 0, 3, 2, 2, 2, 7, 0, 1, 7, 1, 1, 8, 1, 3, 8, 2, 2, 75, 1, 1, 78, 0, 7, 78, 1, 5, 
/* out0432_had-eta12-phi21*/	5, 2, 2, 3, 7, 1, 6, 74, 0, 1, 78, 1, 10, 78, 2, 2, 
/* out0433_had-eta13-phi21*/	7, 1, 0, 6, 7, 1, 3, 74, 0, 2, 74, 2, 3, 77, 0, 1, 77, 1, 3, 78, 2, 1, 
/* out0434_had-eta14-phi21*/	5, 1, 0, 1, 1, 2, 5, 73, 0, 2, 74, 2, 1, 77, 1, 6, 
/* out0435_had-eta15-phi21*/	6, 0, 0, 1, 1, 2, 4, 6, 1, 1, 73, 0, 6, 73, 2, 2, 77, 1, 1, 
/* out0436_had-eta16-phi21*/	2, 0, 0, 5, 73, 2, 6, 
/* out0437_had-eta17-phi21*/	3, 0, 0, 2, 72, 0, 4, 73, 2, 1, 
/* out0438_had-eta18-phi21*/	1, 72, 0, 4, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 132, 0, 2, 
/* out0442_had-eta2-phi22*/	1, 132, 0, 6, 
/* out0443_had-eta3-phi22*/	1, 131, 0, 5, 
/* out0444_had-eta4-phi22*/	1, 131, 0, 3, 
/* out0445_had-eta5-phi22*/	0, 
/* out0446_had-eta6-phi22*/	3, 5, 1, 5, 10, 0, 2, 10, 1, 2, 
/* out0447_had-eta7-phi22*/	3, 4, 0, 8, 5, 1, 4, 10, 1, 12, 
/* out0448_had-eta8-phi22*/	3, 4, 0, 3, 4, 2, 12, 9, 1, 5, 
/* out0449_had-eta9-phi22*/	3, 3, 0, 12, 3, 2, 2, 9, 1, 2, 
/* out0450_had-eta10-phi22*/	3, 2, 0, 2, 3, 2, 11, 8, 1, 1, 
/* out0451_had-eta11-phi22*/	5, 2, 0, 9, 2, 1, 1, 2, 2, 1, 75, 0, 1, 75, 1, 9, 
/* out0452_had-eta12-phi22*/	5, 2, 1, 1, 2, 2, 9, 74, 0, 8, 75, 1, 4, 78, 1, 1, 
/* out0453_had-eta13-phi22*/	6, 1, 0, 7, 1, 1, 1, 2, 2, 1, 74, 0, 4, 74, 1, 2, 74, 2, 5, 
/* out0454_had-eta14-phi22*/	5, 1, 0, 1, 1, 1, 3, 1, 2, 2, 73, 0, 3, 74, 2, 6, 
/* out0455_had-eta15-phi22*/	5, 0, 0, 1, 1, 1, 1, 1, 2, 4, 73, 0, 5, 73, 1, 2, 
/* out0456_had-eta16-phi22*/	4, 0, 0, 3, 0, 1, 4, 73, 1, 3, 73, 2, 4, 
/* out0457_had-eta17-phi22*/	4, 0, 1, 5, 72, 0, 3, 72, 1, 1, 73, 2, 2, 
/* out0458_had-eta18-phi22*/	2, 72, 0, 1, 72, 1, 6, 
/* out0459_had-eta19-phi22*/	1, 72, 1, 1, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 132, 0, 2, 
/* out0462_had-eta2-phi23*/	1, 132, 0, 6, 
/* out0463_had-eta3-phi23*/	1, 131, 0, 5, 
/* out0464_had-eta4-phi23*/	1, 131, 0, 3, 
/* out0465_had-eta5-phi23*/	0, 
/* out0466_had-eta6-phi23*/	2, 5, 0, 9, 5, 1, 2, 
/* out0467_had-eta7-phi23*/	4, 4, 0, 5, 4, 1, 4, 5, 0, 7, 5, 1, 5, 
/* out0468_had-eta8-phi23*/	2, 4, 1, 12, 4, 2, 4, 
/* out0469_had-eta9-phi23*/	2, 3, 0, 3, 3, 1, 9, 
/* out0470_had-eta10-phi23*/	3, 2, 0, 1, 3, 1, 7, 3, 2, 2, 
/* out0471_had-eta11-phi23*/	3, 2, 0, 1, 2, 1, 8, 75, 0, 12, 
/* out0472_had-eta12-phi23*/	5, 2, 1, 6, 74, 0, 1, 74, 1, 2, 75, 0, 3, 75, 1, 2, 
/* out0473_had-eta13-phi23*/	3, 1, 0, 1, 1, 1, 3, 74, 1, 9, 
/* out0474_had-eta14-phi23*/	3, 1, 1, 6, 74, 1, 3, 74, 2, 1, 
/* out0475_had-eta15-phi23*/	2, 1, 1, 2, 73, 1, 5, 
/* out0476_had-eta16-phi23*/	2, 0, 1, 3, 73, 1, 5, 
/* out0477_had-eta17-phi23*/	3, 0, 1, 4, 72, 1, 1, 73, 1, 1, 
/* out0478_had-eta18-phi23*/	1, 72, 1, 5, 
/* out0479_had-eta19-phi23*/	1, 72, 1, 2, 
};