parameter integer matrixH [0:8027] = {
/* num inputs = 152(in0-in151) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 13 */
//* total number of input in adders 2515 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	3,119,1,4,131,0,13,131,1,4,
/* out0004_em-eta4-phi0*/	7,106,1,4,119,1,12,119,2,16,120,0,8,120,1,2,131,0,3,131,2,2,
/* out0005_em-eta5-phi0*/	6,106,1,12,106,2,11,107,0,3,107,1,1,120,0,6,120,2,1,
/* out0006_em-eta6-phi0*/	3,93,1,14,106,2,5,107,0,9,
/* out0007_em-eta7-phi0*/	8,81,1,1,93,1,2,93,2,16,94,0,5,54,0,1,54,1,3,63,1,6,63,2,14,
/* out0008_em-eta8-phi0*/	6,81,1,11,81,2,4,94,0,2,54,0,14,54,1,3,54,2,2,
/* out0009_em-eta9-phi0*/	7,64,1,3,81,2,9,82,0,3,45,0,5,45,1,3,54,0,1,54,2,2,
/* out0010_em-eta10-phi0*/	4,64,1,12,64,2,4,45,0,11,45,2,1,
/* out0011_em-eta11-phi0*/	5,64,2,9,65,0,3,35,0,4,35,1,2,45,2,1,
/* out0012_em-eta12-phi0*/	7,45,4,15,45,5,6,46,0,9,46,1,16,64,2,1,65,0,2,35,0,9,
/* out0013_em-eta13-phi0*/	8,45,5,2,46,0,7,46,4,15,46,5,6,25,0,1,25,1,1,35,0,1,35,2,1,
/* out0014_em-eta14-phi0*/	7,27,4,3,28,1,12,46,2,14,46,3,16,46,4,1,46,5,1,25,0,6,
/* out0015_em-eta15-phi0*/	5,27,4,9,27,5,2,28,0,4,28,1,4,25,0,4,
/* out0016_em-eta16-phi0*/	4,27,5,1,28,0,9,28,4,6,17,2,1,
/* out0017_em-eta17-phi0*/	6,28,2,3,28,3,3,28,4,6,28,5,2,17,0,1,17,2,4,
/* out0018_em-eta18-phi0*/	3,12,3,10,28,2,6,28,3,13,
/* out0019_em-eta19-phi0*/	6,11,0,1,11,1,16,11,2,16,11,3,5,12,3,5,12,4,16,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	6,131,1,12,131,2,8,132,0,3,132,1,2,140,1,3,140,2,13,
/* out0024_em-eta4-phi1*/	6,120,0,1,120,1,14,120,2,3,121,0,1,131,2,6,132,0,11,
/* out0025_em-eta5-phi1*/	4,107,1,10,120,0,1,120,2,12,121,0,6,
/* out0026_em-eta6-phi1*/	5,107,0,4,107,1,5,107,2,15,108,0,1,64,1,1,
/* out0027_em-eta7-phi1*/	8,94,0,5,94,1,13,94,2,2,54,1,3,63,1,10,63,2,2,64,0,12,64,1,1,
/* out0028_em-eta8-phi1*/	10,81,1,4,81,2,3,82,0,1,82,1,4,94,0,4,94,2,8,54,1,7,54,2,9,55,0,3,64,0,2,
/* out0029_em-eta9-phi1*/	6,82,0,8,82,1,4,82,2,1,45,1,11,54,2,3,55,0,5,
/* out0030_em-eta10-phi1*/	9,64,1,1,64,2,1,65,1,2,66,1,7,82,0,4,82,2,4,45,1,2,45,2,12,46,0,1,
/* out0031_em-eta11-phi1*/	8,64,2,1,65,0,6,65,1,14,65,2,9,66,0,2,66,1,4,35,1,10,45,2,1,
/* out0032_em-eta12-phi1*/	9,45,4,1,45,5,4,65,0,5,65,2,4,65,3,15,66,3,3,35,0,2,35,1,1,35,2,7,
/* out0033_em-eta13-phi1*/	8,45,5,4,46,5,9,47,1,8,48,1,2,65,3,1,66,3,2,25,1,5,35,2,3,
/* out0034_em-eta14-phi1*/	8,46,2,2,47,0,12,47,1,6,47,2,1,47,3,1,25,0,3,25,1,3,25,2,1,
/* out0035_em-eta15-phi1*/	6,27,4,4,27,5,5,47,0,4,47,3,7,25,0,2,25,2,4,
/* out0036_em-eta16-phi1*/	6,27,5,8,28,0,3,28,4,4,28,5,7,17,2,5,25,2,1,
/* out0037_em-eta17-phi1*/	6,28,2,4,28,5,6,29,0,2,29,1,1,17,0,3,17,2,3,
/* out0038_em-eta18-phi1*/	4,11,3,2,12,3,1,28,2,3,29,0,6,
/* out0039_em-eta19-phi1*/	3,11,0,4,11,3,9,29,0,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	1,141,1,1,
/* out0043_em-eta3-phi2*/	6,132,1,11,140,1,13,140,2,3,141,0,16,141,1,3,141,2,1,
/* out0044_em-eta4-phi2*/	5,121,1,7,132,0,2,132,1,3,132,2,16,133,0,7,
/* out0045_em-eta5-phi2*/	3,121,0,9,121,1,8,121,2,13,
/* out0046_em-eta6-phi2*/	9,107,2,1,108,0,10,108,1,10,108,2,1,121,2,1,64,1,3,71,0,4,71,1,2,71,2,2,
/* out0047_em-eta7-phi2*/	13,94,1,3,94,2,3,95,0,2,95,1,3,108,0,5,108,2,5,64,0,2,64,1,11,64,2,11,65,0,1,71,0,5,71,1,5,71,2,1,
/* out0048_em-eta8-phi2*/	7,82,1,2,94,2,3,95,0,11,55,0,2,55,1,13,64,2,5,65,0,1,
/* out0049_em-eta9-phi2*/	7,82,1,6,82,2,6,83,0,1,95,0,1,46,1,1,55,0,6,55,2,10,
/* out0050_em-eta10-phi2*/	7,65,4,13,66,1,2,82,2,5,83,0,3,45,2,1,46,0,8,46,1,6,
/* out0051_em-eta11-phi2*/	10,65,2,2,65,4,3,65,5,9,66,0,14,66,1,3,66,4,6,66,5,2,35,1,3,46,0,7,46,2,3,
/* out0052_em-eta12-phi2*/	8,65,2,1,66,2,9,66,3,10,66,4,10,66,5,3,35,2,4,36,0,5,36,1,1,
/* out0053_em-eta13-phi2*/	8,47,1,1,47,4,5,48,0,4,48,1,14,66,3,1,25,1,3,35,2,1,36,0,5,
/* out0054_em-eta14-phi2*/	6,47,1,1,47,2,13,48,0,5,48,4,3,25,1,4,25,2,3,
/* out0055_em-eta15-phi2*/	6,47,2,2,47,3,7,48,3,7,48,4,3,25,2,6,26,0,1,
/* out0056_em-eta16-phi2*/	7,28,5,1,29,1,3,30,1,6,47,3,1,48,3,3,17,0,3,17,2,3,
/* out0057_em-eta17-phi2*/	4,29,1,11,29,2,2,30,1,1,17,0,4,
/* out0058_em-eta18-phi2*/	4,29,0,5,29,1,1,29,2,2,29,3,3,
/* out0059_em-eta19-phi2*/	3,11,0,11,29,0,2,29,3,7,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	4,141,1,3,148,0,9,148,1,3,148,2,6,
/* out0063_em-eta3-phi3*/	8,133,1,3,141,1,9,141,2,15,142,0,10,142,1,2,148,0,6,148,1,11,148,2,7,
/* out0064_em-eta4-phi3*/	4,133,0,8,133,1,13,133,2,13,142,0,1,
/* out0065_em-eta5-phi3*/	7,121,1,1,121,2,2,122,0,11,122,1,10,122,2,2,133,0,1,133,2,2,
/* out0066_em-eta6-phi3*/	8,108,1,6,108,2,5,109,0,3,109,1,2,122,0,5,122,2,3,71,0,1,72,0,4,
/* out0067_em-eta7-phi3*/	11,95,1,9,108,2,5,109,0,7,65,0,6,65,1,13,65,2,1,71,0,6,71,1,9,71,2,13,72,0,3,72,2,1,
/* out0068_em-eta8-phi3*/	8,95,0,2,95,1,4,95,2,11,55,1,3,55,2,1,56,1,3,65,0,8,65,2,7,
/* out0069_em-eta9-phi3*/	7,83,0,2,83,1,8,95,2,3,46,1,1,55,2,5,56,0,11,56,1,1,
/* out0070_em-eta10-phi3*/	6,83,0,9,83,1,1,83,2,2,46,1,8,46,2,4,56,0,2,
/* out0071_em-eta11-phi3*/	9,65,5,7,66,5,8,67,1,7,68,1,4,83,0,1,83,2,2,36,1,3,46,2,9,47,0,1,
/* out0072_em-eta12-phi3*/	9,47,4,1,66,2,7,66,5,3,67,0,13,67,1,8,67,3,1,36,0,2,36,1,8,36,2,1,
/* out0073_em-eta13-phi3*/	7,47,4,10,47,5,10,48,0,2,67,0,3,67,3,2,36,0,4,36,2,5,
/* out0074_em-eta14-phi3*/	8,47,5,2,48,0,5,48,4,8,48,5,7,25,2,1,26,0,2,26,1,3,36,2,1,
/* out0075_em-eta15-phi3*/	5,48,2,11,48,3,5,48,4,2,48,5,1,26,0,6,
/* out0076_em-eta16-phi3*/	5,29,4,6,30,1,8,48,3,1,17,0,2,26,0,3,
/* out0077_em-eta17-phi3*/	4,29,2,3,30,0,9,30,1,1,17,0,3,
/* out0078_em-eta18-phi3*/	3,29,2,8,29,3,1,30,4,3,
/* out0079_em-eta19-phi3*/	4,29,2,1,29,3,5,30,3,4,30,4,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	2,149,0,14,149,1,7,
/* out0083_em-eta3-phi4*/	11,142,0,4,142,1,14,142,2,12,143,0,2,143,2,5,148,0,1,148,1,2,148,2,3,149,0,2,149,1,1,149,2,12,
/* out0084_em-eta4-phi4*/	7,133,2,1,134,0,12,134,1,13,134,2,4,142,0,1,142,2,4,143,2,1,
/* out0085_em-eta5-phi4*/	6,122,1,6,122,2,7,123,0,5,123,1,3,134,0,4,134,2,4,
/* out0086_em-eta6-phi4*/	6,109,1,13,109,2,1,122,2,4,123,0,5,72,0,2,72,1,6,
/* out0087_em-eta7-phi4*/	10,96,1,2,109,0,6,109,2,12,65,1,3,65,2,3,66,0,2,66,1,4,72,0,7,72,1,6,72,2,14,
/* out0088_em-eta8-phi4*/	6,95,2,2,96,0,10,96,1,4,56,1,6,65,2,5,66,0,10,
/* out0089_em-eta9-phi4*/	6,83,1,7,83,2,1,96,0,6,56,0,2,56,1,6,56,2,10,
/* out0090_em-eta10-phi4*/	6,83,2,10,84,0,1,47,0,2,47,1,7,56,0,1,56,2,4,
/* out0091_em-eta11-phi4*/	8,67,4,12,67,5,1,68,0,7,68,1,12,83,2,1,47,0,11,47,1,1,47,2,1,
/* out0092_em-eta12-phi4*/	10,67,1,1,67,2,16,67,3,2,68,0,6,68,4,7,36,1,4,36,2,3,37,0,1,47,0,2,47,2,1,
/* out0093_em-eta13-phi4*/	7,47,5,3,50,1,2,67,3,11,68,3,10,68,4,1,36,2,6,37,0,2,
/* out0094_em-eta14-phi4*/	6,47,5,1,48,2,1,48,5,8,49,1,11,50,1,2,26,1,7,
/* out0095_em-eta15-phi4*/	7,29,4,1,48,2,4,49,0,12,49,1,2,26,0,2,26,1,2,26,2,2,
/* out0096_em-eta16-phi4*/	5,29,4,9,29,5,5,49,0,2,26,0,2,26,2,3,
/* out0097_em-eta17-phi4*/	3,29,5,3,30,0,7,30,4,3,
/* out0098_em-eta18-phi4*/	4,30,2,1,30,3,5,30,4,9,30,5,1,
/* out0099_em-eta19-phi4*/	2,30,2,2,30,3,7,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	1,149,1,5,
/* out0103_em-eta3-phi5*/	5,143,0,14,143,1,11,143,2,6,149,1,3,149,2,4,
/* out0104_em-eta4-phi5*/	6,134,1,3,134,2,6,135,0,9,135,1,8,143,1,5,143,2,4,
/* out0105_em-eta5-phi5*/	5,123,0,2,123,1,13,123,2,6,134,2,2,135,0,7,
/* out0106_em-eta6-phi5*/	9,109,1,1,109,2,1,110,0,1,110,1,7,123,0,4,123,2,10,72,1,1,73,0,1,73,1,2,
/* out0107_em-eta7-phi5*/	11,96,1,3,109,2,2,110,0,14,110,1,1,66,1,11,66,2,1,72,1,3,72,2,1,73,0,15,73,1,4,73,2,8,
/* out0108_em-eta8-phi5*/	7,96,1,7,96,2,9,110,0,1,57,1,3,66,0,4,66,1,1,66,2,15,
/* out0109_em-eta9-phi5*/	6,84,0,1,84,1,6,96,2,7,56,2,2,57,0,10,57,1,5,
/* out0110_em-eta10-phi5*/	5,84,0,10,84,1,2,47,1,8,47,2,1,57,0,6,
/* out0111_em-eta11-phi5*/	6,67,4,4,67,5,15,68,0,1,68,5,3,84,0,4,47,2,12,
/* out0112_em-eta12-phi5*/	8,68,0,2,68,2,8,68,3,1,68,4,8,68,5,13,37,0,2,37,1,8,47,2,1,
/* out0113_em-eta13-phi5*/	5,49,4,8,50,1,5,68,2,8,68,3,5,37,0,8,
/* out0114_em-eta14-phi5*/	7,49,1,2,49,2,5,50,0,8,50,1,7,26,1,4,26,2,1,37,0,3,
/* out0115_em-eta15-phi5*/	5,49,0,1,49,1,1,49,2,11,49,3,5,26,2,6,
/* out0116_em-eta16-phi5*/	4,29,5,4,49,0,1,49,3,11,26,2,4,
/* out0117_em-eta17-phi5*/	2,29,5,4,30,5,9,
/* out0118_em-eta18-phi5*/	2,30,2,5,30,5,6,
/* out0119_em-eta19-phi5*/	1,30,2,8,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	2,150,0,8,150,1,3,
/* out0123_em-eta3-phi6*/	5,144,0,15,144,1,11,144,2,3,150,0,8,150,2,5,
/* out0124_em-eta4-phi6*/	6,135,1,8,135,2,9,136,0,6,136,1,3,144,0,1,144,2,12,
/* out0125_em-eta5-phi6*/	5,124,0,6,124,1,13,124,2,1,135,2,7,136,0,2,
/* out0126_em-eta6-phi6*/	9,110,1,7,110,2,1,111,0,1,111,1,1,124,0,10,124,2,4,73,1,2,74,0,1,74,1,1,
/* out0127_em-eta7-phi6*/	10,97,1,3,110,1,1,110,2,14,111,0,2,67,0,1,67,1,11,73,1,8,73,2,8,74,0,10,74,2,1,
/* out0128_em-eta8-phi6*/	7,97,0,9,97,1,7,110,2,1,57,1,3,67,0,15,67,1,1,67,2,4,
/* out0129_em-eta9-phi6*/	6,84,1,6,84,2,1,97,0,7,57,1,5,57,2,10,58,0,2,
/* out0130_em-eta10-phi6*/	5,84,1,2,84,2,10,48,0,1,48,1,8,57,2,6,
/* out0131_em-eta11-phi6*/	6,69,1,3,69,4,4,70,0,1,70,1,15,84,2,4,48,0,12,
/* out0132_em-eta12-phi6*/	8,69,0,8,69,1,13,69,2,8,69,3,1,70,0,2,37,1,8,37,2,2,48,0,1,
/* out0133_em-eta13-phi6*/	5,49,4,8,49,5,5,69,0,8,69,3,5,37,2,8,
/* out0134_em-eta14-phi6*/	7,49,5,7,50,0,8,50,4,5,50,5,2,27,0,1,27,1,4,37,2,3,
/* out0135_em-eta15-phi6*/	5,50,2,1,50,3,5,50,4,11,50,5,1,27,0,6,
/* out0136_em-eta16-phi6*/	4,32,1,4,50,2,1,50,3,11,27,0,4,
/* out0137_em-eta17-phi6*/	2,31,1,9,32,1,4,
/* out0138_em-eta18-phi6*/	2,31,0,5,31,1,6,
/* out0139_em-eta19-phi6*/	1,31,0,8,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	1,150,1,11,
/* out0143_em-eta3-phi7*/	9,144,1,5,145,0,12,145,1,14,145,2,4,150,1,2,150,2,11,151,0,3,151,1,2,151,2,1,
/* out0144_em-eta4-phi7*/	7,136,0,4,136,1,13,136,2,12,137,0,1,144,2,1,145,0,4,145,2,1,
/* out0145_em-eta5-phi7*/	6,124,1,3,124,2,5,125,0,7,125,1,6,136,0,4,136,2,4,
/* out0146_em-eta6-phi7*/	5,111,0,1,111,1,13,124,2,6,125,0,4,74,1,7,
/* out0147_em-eta7-phi7*/	10,97,1,2,111,0,12,111,2,6,67,1,4,67,2,2,68,0,3,68,1,3,74,0,5,74,1,6,74,2,14,
/* out0148_em-eta8-phi7*/	6,97,1,4,97,2,10,98,0,2,58,1,6,67,2,10,68,0,5,
/* out0149_em-eta9-phi7*/	6,85,0,1,85,1,7,97,2,6,58,0,10,58,1,6,58,2,2,
/* out0150_em-eta10-phi7*/	6,84,2,1,85,0,10,48,1,7,48,2,2,58,0,4,58,2,1,
/* out0151_em-eta11-phi7*/	8,69,4,12,69,5,12,70,0,7,70,1,1,85,0,1,48,0,1,48,1,1,48,2,11,
/* out0152_em-eta12-phi7*/	10,69,2,7,70,0,6,70,3,2,70,4,16,70,5,1,37,2,1,38,0,3,38,1,4,48,0,1,48,2,2,
/* out0153_em-eta13-phi7*/	7,49,5,2,52,1,3,69,2,1,69,3,10,70,3,11,37,2,2,38,0,6,
/* out0154_em-eta14-phi7*/	6,49,5,2,50,5,11,51,0,1,51,1,8,52,1,1,27,1,7,
/* out0155_em-eta15-phi7*/	7,31,4,1,50,2,12,50,5,2,51,0,4,27,0,2,27,1,2,27,2,2,
/* out0156_em-eta16-phi7*/	5,31,4,9,32,1,5,50,2,2,27,0,3,27,2,2,
/* out0157_em-eta17-phi7*/	3,31,2,3,32,0,7,32,1,3,
/* out0158_em-eta18-phi7*/	4,31,0,1,31,1,1,31,2,9,31,3,5,
/* out0159_em-eta19-phi7*/	2,31,0,2,31,3,7,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	4,146,1,3,151,0,6,151,1,3,151,2,9,
/* out0163_em-eta3-phi8*/	8,137,1,3,145,1,2,145,2,10,146,0,15,146,1,9,151,0,7,151,1,11,151,2,6,
/* out0164_em-eta4-phi8*/	4,137,0,13,137,1,13,137,2,8,145,2,1,
/* out0165_em-eta5-phi8*/	7,125,0,2,125,1,10,125,2,11,126,0,2,126,1,1,137,0,2,137,2,1,
/* out0166_em-eta6-phi8*/	8,111,1,2,111,2,3,112,0,5,112,1,6,125,0,3,125,2,5,74,1,1,75,2,1,
/* out0167_em-eta7-phi8*/	11,98,1,9,111,2,7,112,0,5,68,0,1,68,1,13,68,2,6,74,1,1,74,2,1,75,0,13,75,1,9,75,2,6,
/* out0168_em-eta8-phi8*/	8,98,0,11,98,1,4,98,2,2,58,1,3,59,0,1,59,1,3,68,0,7,68,2,8,
/* out0169_em-eta9-phi8*/	7,85,1,8,85,2,2,98,0,3,49,1,1,58,1,1,58,2,11,59,0,5,
/* out0170_em-eta10-phi8*/	6,85,0,2,85,1,1,85,2,9,49,0,4,49,1,8,58,2,2,
/* out0171_em-eta11-phi8*/	9,69,5,4,70,5,7,71,1,8,72,1,7,85,0,2,85,2,1,38,1,3,48,2,1,49,0,9,
/* out0172_em-eta12-phi8*/	9,51,4,1,70,2,13,70,3,1,70,5,8,71,0,7,71,1,3,38,0,1,38,1,8,38,2,2,
/* out0173_em-eta13-phi8*/	7,51,4,10,52,0,2,52,1,10,70,2,3,70,3,2,38,0,5,38,2,4,
/* out0174_em-eta14-phi8*/	8,51,1,7,51,2,8,52,0,5,52,1,2,27,1,3,27,2,2,28,0,1,38,0,1,
/* out0175_em-eta15-phi8*/	5,51,0,11,51,1,1,51,2,2,51,3,5,27,2,6,
/* out0176_em-eta16-phi8*/	5,31,4,6,31,5,8,51,3,1,18,1,2,27,2,3,
/* out0177_em-eta17-phi8*/	4,31,5,1,32,0,9,32,4,3,18,1,3,
/* out0178_em-eta18-phi8*/	3,31,2,3,32,3,1,32,4,8,
/* out0179_em-eta19-phi8*/	4,31,2,1,31,3,4,32,3,5,32,4,1,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	1,146,1,1,
/* out0183_em-eta3-phi9*/	6,138,1,11,146,0,1,146,1,3,146,2,16,147,0,12,147,2,4,
/* out0184_em-eta4-phi9*/	5,126,1,7,137,2,7,138,0,16,138,1,3,138,2,2,
/* out0185_em-eta5-phi9*/	3,126,0,13,126,1,8,126,2,9,
/* out0186_em-eta6-phi9*/	9,112,0,1,112,1,10,112,2,10,113,0,1,126,0,1,69,1,3,75,0,2,75,1,2,75,2,4,
/* out0187_em-eta7-phi9*/	13,98,1,3,98,2,2,99,0,3,99,1,3,112,0,5,112,2,5,68,2,1,69,0,11,69,1,11,69,2,2,75,0,1,75,1,5,75,2,5,
/* out0188_em-eta8-phi9*/	7,86,1,2,98,2,11,99,0,3,59,1,13,59,2,2,68,2,1,69,0,5,
/* out0189_em-eta9-phi9*/	7,85,2,1,86,0,6,86,1,6,98,2,1,49,1,1,59,0,10,59,2,6,
/* out0190_em-eta10-phi9*/	7,71,4,13,71,5,2,85,2,3,86,0,5,49,1,6,49,2,8,50,0,1,
/* out0191_em-eta11-phi9*/	10,71,1,2,71,2,6,71,4,3,71,5,3,72,0,14,72,1,9,72,4,2,39,1,3,49,0,3,49,2,7,
/* out0192_em-eta12-phi9*/	8,71,0,9,71,1,3,71,2,10,71,3,10,72,4,1,38,1,1,38,2,5,39,0,4,
/* out0193_em-eta13-phi9*/	8,51,4,5,51,5,14,52,0,4,52,5,1,71,3,1,28,1,3,38,2,5,39,0,1,
/* out0194_em-eta14-phi9*/	6,51,2,3,52,0,5,52,4,13,52,5,1,28,0,3,28,1,4,
/* out0195_em-eta15-phi9*/	6,51,2,3,51,3,7,52,3,7,52,4,2,27,2,1,28,0,6,
/* out0196_em-eta16-phi9*/	7,31,5,6,32,5,3,33,1,1,51,3,3,52,3,1,18,1,3,18,2,3,
/* out0197_em-eta17-phi9*/	4,31,5,1,32,4,2,32,5,11,18,1,4,
/* out0198_em-eta18-phi9*/	4,32,2,5,32,3,3,32,4,2,32,5,1,
/* out0199_em-eta19-phi9*/	3,13,4,11,32,2,2,32,3,7,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	6,138,1,2,138,2,3,139,0,8,139,1,12,147,0,4,147,2,12,
/* out0204_em-eta4-phi10*/	6,126,2,1,127,0,3,127,1,14,127,2,1,138,2,11,139,0,6,
/* out0205_em-eta5-phi10*/	4,113,1,10,126,2,6,127,0,12,127,2,1,
/* out0206_em-eta6-phi10*/	6,112,2,1,113,0,15,113,1,5,113,2,4,69,1,1,70,0,1,
/* out0207_em-eta7-phi10*/	8,99,0,2,99,1,13,99,2,5,60,1,3,69,1,1,69,2,12,70,0,10,70,2,2,
/* out0208_em-eta8-phi10*/	8,86,1,4,86,2,1,99,0,8,99,2,4,59,2,3,60,0,9,60,1,7,69,2,2,
/* out0209_em-eta9-phi10*/	6,86,0,1,86,1,4,86,2,8,50,1,11,59,2,5,60,0,3,
/* out0210_em-eta10-phi10*/	9,71,5,7,72,5,2,73,0,1,73,1,1,86,0,4,86,2,4,49,2,1,50,0,12,50,1,2,
/* out0211_em-eta11-phi10*/	7,71,5,4,72,0,2,72,2,6,72,4,9,72,5,14,39,1,10,50,0,1,
/* out0212_em-eta12-phi10*/	9,53,4,1,54,1,4,71,3,3,72,2,5,72,3,15,72,4,4,39,0,7,39,1,1,39,2,2,
/* out0213_em-eta13-phi10*/	8,51,5,2,52,5,8,53,1,9,54,1,4,71,3,2,72,3,1,28,1,5,39,0,3,
/* out0214_em-eta14-phi10*/	8,52,2,12,52,3,1,52,4,1,52,5,6,53,0,2,28,0,1,28,1,3,28,2,3,
/* out0215_em-eta15-phi10*/	6,33,4,4,34,1,5,52,2,4,52,3,7,28,0,4,28,2,2,
/* out0216_em-eta16-phi10*/	4,33,1,7,34,1,8,18,2,5,28,0,1,
/* out0217_em-eta17-phi10*/	6,32,2,2,32,5,1,33,0,4,33,1,6,18,1,3,18,2,3,
/* out0218_em-eta18-phi10*/	4,13,5,2,14,5,1,32,2,6,33,0,3,
/* out0219_em-eta19-phi10*/	3,13,4,4,13,5,9,32,2,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	2,139,1,4,139,2,13,
/* out0224_em-eta4-phi11*/	5,127,1,2,127,2,8,128,2,5,139,0,2,139,2,3,
/* out0225_em-eta5-phi11*/	6,113,1,1,113,2,3,114,0,7,114,1,12,127,0,1,127,2,6,
/* out0226_em-eta6-phi11*/	3,100,1,10,113,2,9,114,0,5,
/* out0227_em-eta7-phi11*/	10,87,1,1,99,2,5,100,0,12,100,1,2,60,1,3,60,2,1,61,0,2,61,1,4,70,0,5,70,2,14,
/* out0228_em-eta8-phi11*/	8,87,0,3,87,1,11,99,2,2,51,1,1,60,0,2,60,1,3,60,2,14,61,0,2,
/* out0229_em-eta9-phi11*/	9,73,1,2,86,2,3,87,0,9,50,1,3,50,2,5,51,0,4,51,1,3,60,0,2,60,2,1,
/* out0230_em-eta10-phi11*/	5,73,0,2,73,1,9,40,1,3,50,0,1,50,2,11,
/* out0231_em-eta11-phi11*/	7,72,2,3,73,0,9,39,1,2,39,2,5,40,0,4,40,1,1,50,0,1,
/* out0232_em-eta12-phi11*/	7,53,4,15,53,5,4,54,0,5,54,1,6,72,2,2,29,1,2,39,2,8,
/* out0233_em-eta13-phi11*/	10,53,1,6,53,2,11,54,0,7,54,1,2,28,1,1,28,2,1,29,0,3,29,1,2,39,0,1,39,2,1,
/* out0234_em-eta14-phi11*/	7,33,4,3,53,0,14,53,1,1,53,2,1,53,3,4,28,2,6,29,0,1,
/* out0235_em-eta15-phi11*/	6,33,4,9,33,5,4,34,0,3,34,1,2,19,1,3,28,2,4,
/* out0236_em-eta16-phi11*/	6,33,2,6,34,0,9,34,1,1,18,2,1,19,0,3,19,1,1,
/* out0237_em-eta17-phi11*/	7,33,0,3,33,1,2,33,2,6,33,3,3,18,1,1,18,2,4,19,0,1,
/* out0238_em-eta18-phi11*/	3,14,5,6,33,0,6,33,3,1,
/* out0239_em-eta19-phi11*/	6,13,4,1,13,5,5,14,0,15,14,1,16,14,4,4,14,5,5,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	4,128,1,1,128,2,1,129,0,6,129,1,12,
/* out0244_em-eta4-phi12*/	5,115,0,1,115,1,9,128,1,15,128,2,10,129,0,5,
/* out0245_em-eta5-phi12*/	5,101,1,3,114,0,1,114,1,4,114,2,14,115,0,7,
/* out0246_em-eta6-phi12*/	6,100,1,4,100,2,7,101,0,6,101,1,4,114,0,3,114,2,2,
/* out0247_em-eta7-phi12*/	9,87,1,1,88,0,1,88,1,4,100,0,4,100,2,9,61,0,3,61,1,12,61,2,9,62,0,1,
/* out0248_em-eta8-phi12*/	7,87,1,3,87,2,11,88,0,2,51,1,8,51,2,2,61,0,9,61,2,2,
/* out0249_em-eta9-phi12*/	9,73,1,2,73,2,1,74,0,1,74,1,2,87,0,4,87,2,5,51,0,8,51,1,4,51,2,6,
/* out0250_em-eta10-phi12*/	5,73,1,2,73,2,9,40,1,10,40,2,1,51,0,4,
/* out0251_em-eta11-phi12*/	6,56,1,3,73,0,4,73,2,5,40,0,8,40,1,2,40,2,2,
/* out0252_em-eta12-phi12*/	7,53,5,12,54,0,3,54,4,2,54,5,13,55,1,2,29,1,7,40,0,3,
/* out0253_em-eta13-phi12*/	9,53,2,3,54,0,1,54,2,1,54,3,6,54,4,14,54,5,2,29,0,4,29,1,4,29,2,1,
/* out0254_em-eta14-phi12*/	6,33,5,3,53,2,1,53,3,12,54,3,6,19,1,1,29,0,6,
/* out0255_em-eta15-phi12*/	5,33,5,9,34,0,2,34,4,1,34,5,6,19,1,6,
/* out0256_em-eta16-phi12*/	6,33,2,1,34,0,2,34,4,12,34,5,1,19,0,4,19,1,2,
/* out0257_em-eta17-phi12*/	5,33,2,3,33,3,4,34,3,3,34,4,3,19,0,4,
/* out0258_em-eta18-phi12*/	3,14,2,5,14,5,1,33,3,7,
/* out0259_em-eta19-phi12*/	5,14,0,1,14,2,3,14,3,5,14,4,11,14,5,3,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	6,116,1,5,129,0,1,129,1,4,129,2,14,130,0,13,130,2,3,
/* out0264_em-eta4-phi13*/	6,115,1,7,115,2,11,116,0,7,116,1,4,129,0,4,129,2,2,
/* out0265_em-eta5-phi13*/	6,101,1,6,101,2,4,102,0,3,102,1,4,115,0,8,115,2,5,
/* out0266_em-eta6-phi13*/	4,101,0,10,101,1,3,101,2,10,62,0,2,
/* out0267_em-eta7-phi13*/	7,88,0,2,88,1,12,88,2,6,52,1,7,61,2,4,62,0,12,62,2,9,
/* out0268_em-eta8-phi13*/	8,74,1,4,88,0,11,88,2,1,51,2,1,52,0,10,52,1,8,52,2,1,61,2,1,
/* out0269_em-eta9-phi13*/	6,74,0,4,74,1,9,74,2,1,41,1,9,51,2,7,52,0,3,
/* out0270_em-eta10-phi13*/	7,55,4,8,55,5,2,73,2,1,74,0,8,40,2,5,41,0,8,41,1,2,
/* out0271_em-eta11-phi13*/	8,55,1,1,55,2,2,55,4,8,55,5,2,56,0,9,56,1,13,30,1,5,40,2,8,
/* out0272_em-eta12-phi13*/	10,54,2,3,54,5,1,55,0,10,55,1,13,55,2,5,29,1,1,29,2,4,30,0,3,30,1,1,40,0,1,
/* out0273_em-eta13-phi13*/	6,35,4,10,36,1,1,54,2,12,54,3,2,55,0,3,29,2,8,
/* out0274_em-eta14-phi13*/	9,35,1,5,36,1,14,54,3,2,19,1,1,19,2,1,20,0,1,20,1,1,29,0,2,29,2,2,
/* out0275_em-eta15-phi13*/	6,34,2,2,34,5,7,35,0,3,35,1,8,19,1,2,19,2,4,
/* out0276_em-eta16-phi13*/	5,34,2,11,34,3,2,34,5,2,19,0,1,19,2,4,
/* out0277_em-eta17-phi13*/	6,15,4,1,16,1,2,34,2,2,34,3,9,19,0,3,19,2,1,
/* out0278_em-eta18-phi13*/	5,14,2,3,15,1,3,16,1,4,33,3,1,34,3,2,
/* out0279_em-eta19-phi13*/	4,14,2,5,14,3,9,14,4,1,15,1,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	1,117,1,2,
/* out0283_em-eta3-phi14*/	6,116,1,5,116,2,6,117,0,9,117,1,11,130,0,3,130,2,13,
/* out0284_em-eta4-phi14*/	7,102,1,5,102,2,2,103,0,2,103,1,5,116,0,9,116,1,2,116,2,10,
/* out0285_em-eta5-phi14*/	3,102,0,12,102,1,7,102,2,11,
/* out0286_em-eta6-phi14*/	9,89,0,3,89,1,16,89,2,3,101,2,2,102,0,1,53,0,2,53,1,1,62,0,1,62,2,1,
/* out0287_em-eta7-phi14*/	9,75,1,4,88,2,6,89,0,10,52,1,1,52,2,3,53,0,14,53,1,3,53,2,9,62,2,6,
/* out0288_em-eta8-phi14*/	9,74,1,1,74,2,2,75,0,5,75,1,6,88,2,3,42,1,6,52,0,2,52,2,12,53,2,1,
/* out0289_em-eta9-phi14*/	7,57,1,1,74,2,11,75,0,2,41,1,5,41,2,8,42,0,3,52,0,1,
/* out0290_em-eta10-phi14*/	9,55,5,9,56,5,6,57,0,1,57,1,2,74,0,3,74,2,2,30,1,1,41,0,8,41,2,6,
/* out0291_em-eta11-phi14*/	9,55,2,2,55,5,3,56,0,7,56,2,1,56,3,2,56,4,14,56,5,10,30,1,9,30,2,3,
/* out0292_em-eta12-phi14*/	7,55,0,2,55,2,7,55,3,15,56,3,5,56,4,2,30,0,9,30,2,1,
/* out0293_em-eta13-phi14*/	7,35,4,6,35,5,13,36,0,5,55,0,1,20,1,6,29,2,1,30,0,2,
/* out0294_em-eta14-phi14*/	6,35,2,8,36,0,11,36,1,1,36,4,2,20,0,3,20,1,4,
/* out0295_em-eta15-phi14*/	6,35,0,8,35,1,3,35,2,5,35,3,3,19,2,2,20,0,4,
/* out0296_em-eta16-phi14*/	5,15,4,10,34,2,1,35,0,5,11,1,2,19,2,3,
/* out0297_em-eta17-phi14*/	5,15,4,4,16,0,2,16,1,7,11,1,2,19,2,1,
/* out0298_em-eta18-phi14*/	4,15,1,5,15,2,1,16,0,1,16,1,3,
/* out0299_em-eta19-phi14*/	3,14,3,2,15,0,3,15,1,5,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	5,117,1,1,117,2,1,118,0,9,118,1,3,118,2,6,
/* out0303_em-eta3-phi15*/	10,103,1,2,103,2,1,104,0,3,104,1,9,117,0,7,117,1,2,117,2,15,118,0,6,118,1,11,118,2,7,
/* out0304_em-eta4-phi15*/	4,103,0,11,103,1,9,103,2,14,104,0,1,
/* out0305_em-eta5-phi15*/	5,90,0,5,90,1,16,90,2,3,102,2,3,103,0,3,
/* out0306_em-eta6-phi15*/	3,76,1,5,89,2,11,90,0,8,
/* out0307_em-eta7-phi15*/	10,75,1,4,75,2,5,76,0,4,76,1,3,89,0,3,89,2,2,43,0,1,43,1,5,53,1,12,53,2,5,
/* out0308_em-eta8-phi15*/	8,75,0,6,75,1,2,75,2,9,42,0,1,42,1,10,42,2,9,43,0,1,53,2,1,
/* out0309_em-eta9-phi15*/	7,57,1,10,57,2,1,75,0,3,31,1,5,41,2,1,42,0,11,42,2,1,
/* out0310_em-eta10-phi15*/	5,57,0,8,57,1,3,31,0,5,31,1,9,41,2,1,
/* out0311_em-eta11-phi15*/	7,37,4,11,56,2,14,56,3,1,57,0,3,21,1,1,30,2,7,31,0,4,
/* out0312_em-eta12-phi15*/	11,35,5,1,37,1,5,37,4,1,38,1,15,55,3,1,56,2,1,56,3,8,21,0,1,21,1,3,30,0,2,30,2,5,
/* out0313_em-eta13-phi15*/	8,35,5,2,36,2,3,36,4,2,36,5,15,37,0,1,37,1,5,20,1,4,20,2,5,
/* out0314_em-eta14-phi15*/	8,35,2,1,36,2,3,36,3,6,36,4,12,36,5,1,20,0,2,20,1,1,20,2,4,
/* out0315_em-eta15-phi15*/	5,35,2,2,35,3,12,36,3,4,11,2,1,20,0,5,
/* out0316_em-eta16-phi15*/	5,15,4,1,15,5,13,35,3,1,11,1,2,11,2,3,
/* out0317_em-eta17-phi15*/	4,15,5,1,16,0,11,16,4,1,11,1,4,
/* out0318_em-eta18-phi15*/	3,15,2,9,16,0,2,11,1,1,
/* out0319_em-eta19-phi15*/	4,15,0,5,15,1,2,15,2,2,15,3,1,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	1,105,1,12,
/* out0323_em-eta3-phi16*/	11,92,0,2,92,2,5,104,0,7,104,1,7,104,2,16,105,0,16,105,1,1,105,2,5,118,0,1,118,1,2,118,2,3,
/* out0324_em-eta4-phi16*/	6,91,0,6,91,1,16,91,2,7,92,2,1,103,2,1,104,0,5,
/* out0325_em-eta5-phi16*/	3,77,1,8,90,2,12,91,0,9,
/* out0326_em-eta6-phi16*/	11,76,1,7,76,2,8,77,0,4,77,1,2,90,0,3,90,2,1,43,1,1,43,2,1,44,0,3,44,1,2,44,2,1,
/* out0327_em-eta7-phi16*/	9,58,1,2,76,0,12,76,1,1,76,2,4,43,0,5,43,1,10,43,2,10,44,0,1,44,1,1,
/* out0328_em-eta8-phi16*/	6,58,0,2,58,1,12,75,2,2,32,1,9,42,2,4,43,0,9,
/* out0329_em-eta9-phi16*/	8,57,2,8,58,0,6,31,1,1,31,2,4,32,0,6,32,1,4,42,0,1,42,2,2,
/* out0330_em-eta10-phi16*/	6,39,1,1,57,0,3,57,2,7,31,0,2,31,1,1,31,2,12,
/* out0331_em-eta11-phi16*/	9,37,4,4,37,5,16,38,0,5,38,4,2,38,5,6,57,0,1,21,1,7,21,2,1,31,0,5,
/* out0332_em-eta12-phi16*/	8,37,1,2,37,2,13,38,0,11,38,1,1,38,4,5,21,0,4,21,1,5,21,2,1,
/* out0333_em-eta13-phi16*/	9,17,4,2,36,2,3,37,0,14,37,1,4,37,2,1,37,3,3,12,1,1,20,2,2,21,0,6,
/* out0334_em-eta14-phi16*/	6,17,4,9,18,1,4,36,2,7,36,3,2,12,1,3,20,2,4,
/* out0335_em-eta15-phi16*/	9,16,5,1,17,1,4,18,1,9,36,3,4,11,2,3,12,0,1,12,1,1,20,0,1,20,2,1,
/* out0336_em-eta16-phi16*/	4,15,5,2,16,5,12,17,1,2,11,2,6,
/* out0337_em-eta17-phi16*/	4,16,4,10,16,5,3,11,0,2,11,1,3,
/* out0338_em-eta18-phi16*/	5,15,2,4,15,3,1,16,3,1,16,4,5,11,1,1,
/* out0339_em-eta19-phi16*/	2,15,0,8,15,3,9,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	2,105,1,3,105,2,4,
/* out0343_em-eta3-phi17*/	4,92,0,14,92,1,11,92,2,6,105,2,7,
/* out0344_em-eta4-phi17*/	5,78,0,2,78,1,16,91,2,8,92,1,5,92,2,4,
/* out0345_em-eta5-phi17*/	5,77,1,6,77,2,14,78,0,6,91,0,1,91,2,1,
/* out0346_em-eta6-phi17*/	7,59,1,9,76,2,2,77,0,12,77,2,2,44,0,6,44,1,1,44,2,7,
/* out0347_em-eta7-phi17*/	11,58,1,1,58,2,2,59,0,8,59,1,7,76,2,2,33,0,1,33,1,15,43,2,5,44,0,6,44,1,12,44,2,8,
/* out0348_em-eta8-phi17*/	7,58,0,2,58,1,1,58,2,13,32,1,3,32,2,10,33,0,7,33,1,1,
/* out0349_em-eta9-phi17*/	6,39,1,7,58,0,6,58,2,1,22,1,3,32,0,10,32,2,6,
/* out0350_em-eta10-phi17*/	4,39,0,4,39,1,8,22,0,1,22,1,13,
/* out0351_em-eta11-phi17*/	6,38,2,11,38,4,1,38,5,10,39,0,4,21,2,5,22,0,7,
/* out0352_em-eta12-phi17*/	7,37,2,2,37,3,2,38,2,5,38,3,15,38,4,8,21,0,1,21,2,9,
/* out0353_em-eta13-phi17*/	7,17,4,2,17,5,11,37,0,1,37,3,11,38,3,1,12,1,5,21,0,4,
/* out0354_em-eta14-phi17*/	6,17,4,3,17,5,5,18,0,13,18,1,2,12,0,1,12,1,6,
/* out0355_em-eta15-phi17*/	5,17,1,6,17,2,8,18,0,3,18,1,1,12,0,5,
/* out0356_em-eta16-phi17*/	6,16,2,4,17,0,8,17,1,4,11,0,3,11,2,3,12,0,1,
/* out0357_em-eta17-phi17*/	3,16,2,12,16,3,2,11,0,10,
/* out0358_em-eta18-phi17*/	3,16,3,10,11,0,1,11,1,1,
/* out0359_em-eta19-phi17*/	2,15,3,5,16,3,3,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	1,80,1,7,
/* out0363_em-eta3-phi18*/	5,79,0,3,79,1,15,79,2,5,80,0,11,80,1,3,
/* out0364_em-eta4-phi18*/	5,61,1,8,78,0,2,78,2,16,79,0,13,79,2,5,
/* out0365_em-eta5-phi18*/	5,60,1,14,60,2,6,61,0,1,61,1,1,78,0,6,
/* out0366_em-eta6-phi18*/	7,41,1,2,59,2,9,60,0,12,60,1,2,34,0,7,34,1,1,34,2,6,
/* out0367_em-eta7-phi18*/	11,40,1,2,40,2,1,41,1,2,59,0,8,59,2,7,24,1,5,33,0,1,33,2,15,34,0,8,34,1,12,34,2,6,
/* out0368_em-eta8-phi18*/	7,40,0,2,40,1,13,40,2,1,23,1,10,23,2,3,33,0,7,33,2,1,
/* out0369_em-eta9-phi18*/	6,39,2,7,40,0,6,40,1,1,22,2,3,23,0,10,23,1,6,
/* out0370_em-eta10-phi18*/	4,39,0,4,39,2,8,22,0,1,22,2,13,
/* out0371_em-eta11-phi18*/	6,19,4,11,19,5,10,20,0,1,39,0,4,13,1,5,22,0,7,
/* out0372_em-eta12-phi18*/	7,19,1,2,19,2,2,19,4,5,20,0,8,20,1,15,13,0,1,13,1,9,
/* out0373_em-eta13-phi18*/	7,18,2,2,18,5,11,19,0,1,19,1,11,20,1,1,12,2,5,13,0,4,
/* out0374_em-eta14-phi18*/	6,18,2,3,18,3,2,18,4,13,18,5,5,12,0,1,12,2,6,
/* out0375_em-eta15-phi18*/	5,17,2,8,17,3,6,18,3,1,18,4,3,12,0,5,
/* out0376_em-eta16-phi18*/	6,0,4,4,17,0,8,17,3,4,5,1,1,5,2,3,12,0,1,
/* out0377_em-eta17-phi18*/	3,0,4,12,1,1,2,5,1,4,
/* out0378_em-eta18-phi18*/	2,1,1,10,5,1,2,
/* out0379_em-eta19-phi18*/	2,0,1,5,1,1,3,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	2,80,1,6,80,2,6,
/* out0383_em-eta3-phi19*/	10,62,0,7,62,1,16,62,2,7,63,0,3,63,1,2,63,2,1,79,1,1,79,2,5,80,0,5,80,2,10,
/* out0384_em-eta4-phi19*/	6,43,1,1,61,0,6,61,1,7,61,2,16,62,0,5,79,2,1,
/* out0385_em-eta5-phi19*/	3,42,1,12,60,2,8,61,0,9,
/* out0386_em-eta6-phi19*/	11,41,1,8,41,2,7,42,0,3,42,1,1,60,0,4,60,2,2,24,1,1,24,2,1,34,0,1,34,1,2,34,2,3,
/* out0387_em-eta7-phi19*/	9,40,2,2,41,0,12,41,1,4,41,2,1,24,0,5,24,1,10,24,2,10,34,1,1,34,2,1,
/* out0388_em-eta8-phi19*/	6,22,1,2,40,0,2,40,2,12,15,1,4,23,2,9,24,0,9,
/* out0389_em-eta9-phi19*/	8,21,1,8,40,0,6,14,1,4,14,2,1,15,0,1,15,1,2,23,0,6,23,2,4,
/* out0390_em-eta10-phi19*/	6,21,0,3,21,1,7,39,2,1,14,0,2,14,1,12,14,2,1,
/* out0391_em-eta11-phi19*/	9,19,5,6,20,0,2,20,2,4,20,4,5,20,5,16,21,0,1,13,1,1,13,2,7,14,0,5,
/* out0392_em-eta12-phi19*/	8,19,2,13,19,3,2,20,0,5,20,3,1,20,4,11,13,0,4,13,1,1,13,2,5,
/* out0393_em-eta13-phi19*/	9,2,4,3,18,2,2,19,0,14,19,1,3,19,2,1,19,3,4,6,1,2,12,2,1,13,0,6,
/* out0394_em-eta14-phi19*/	6,2,4,7,3,1,2,18,2,9,18,3,4,6,1,4,12,2,3,
/* out0395_em-eta15-phi19*/	9,0,5,1,3,1,4,17,3,4,18,3,9,5,2,3,6,0,1,6,1,1,12,0,1,12,2,1,
/* out0396_em-eta16-phi19*/	4,0,5,12,1,5,2,17,3,2,5,2,5,
/* out0397_em-eta17-phi19*/	3,0,5,3,1,0,10,5,1,4,
/* out0398_em-eta18-phi19*/	5,0,1,1,0,2,4,1,0,5,1,1,1,5,1,1,
/* out0399_em-eta19-phi19*/	2,0,0,8,0,1,9,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	5,44,1,1,44,2,1,63,0,6,63,1,3,63,2,9,
/* out0403_em-eta3-phi20*/	10,43,1,1,43,2,2,44,0,7,44,1,15,44,2,2,62,0,3,62,2,9,63,0,7,63,1,11,63,2,6,
/* out0404_em-eta4-phi20*/	4,43,0,11,43,1,14,43,2,9,62,0,1,
/* out0405_em-eta5-phi20*/	5,24,1,3,42,0,5,42,1,3,42,2,16,43,0,3,
/* out0406_em-eta6-phi20*/	3,23,1,11,41,2,5,42,0,8,
/* out0407_em-eta7-phi20*/	11,22,1,5,22,2,4,23,0,3,23,1,2,41,0,4,41,2,3,16,0,16,16,1,5,16,2,6,24,0,1,24,2,5,
/* out0408_em-eta8-phi20*/	8,22,0,6,22,1,9,22,2,2,15,0,1,15,1,9,15,2,10,16,2,1,24,0,1,
/* out0409_em-eta9-phi20*/	7,21,1,1,21,2,10,22,0,3,8,1,1,14,2,5,15,0,11,15,1,1,
/* out0410_em-eta10-phi20*/	5,21,0,8,21,2,3,8,1,1,14,0,5,14,2,9,
/* out0411_em-eta11-phi20*/	7,4,4,14,5,1,1,20,2,11,21,0,3,7,1,7,13,2,1,14,0,4,
/* out0412_em-eta12-phi20*/	11,3,5,1,4,1,1,4,4,1,5,1,8,19,3,5,20,2,1,20,3,15,7,0,2,7,1,5,13,0,1,13,2,3,
/* out0413_em-eta13-phi20*/	8,2,4,3,2,5,15,3,0,2,3,5,2,19,0,1,19,3,5,6,1,5,6,2,4,
/* out0414_em-eta14-phi20*/	8,2,2,1,2,4,3,2,5,1,3,0,12,3,1,6,6,0,2,6,1,4,6,2,1,
/* out0415_em-eta15-phi20*/	5,2,1,12,2,2,2,3,1,4,5,2,1,6,0,5,
/* out0416_em-eta16-phi20*/	5,1,2,1,1,5,13,2,1,1,5,0,4,5,2,4,
/* out0417_em-eta17-phi20*/	5,1,0,1,1,4,11,1,5,1,5,0,3,5,1,2,
/* out0418_em-eta18-phi20*/	3,0,2,9,1,4,2,5,1,1,
/* out0419_em-eta19-phi20*/	4,0,0,5,0,1,1,0,2,2,0,3,2,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	1,44,2,2,
/* out0423_em-eta3-phi21*/	6,25,1,6,25,2,5,26,0,12,26,2,4,44,0,9,44,2,11,
/* out0424_em-eta4-phi21*/	7,24,1,2,24,2,5,25,0,9,25,1,10,25,2,2,43,0,2,43,2,5,
/* out0425_em-eta5-phi21*/	3,24,0,12,24,1,11,24,2,7,
/* out0426_em-eta6-phi21*/	7,8,1,2,23,0,3,23,1,3,23,2,16,24,0,1,10,0,3,16,1,2,
/* out0427_em-eta7-phi21*/	8,7,1,6,22,2,4,23,0,10,9,1,3,9,2,1,10,0,5,16,1,9,16,2,8,
/* out0428_em-eta8-phi21*/	9,6,1,2,6,2,1,7,1,3,22,0,5,22,2,6,9,0,2,9,1,12,15,2,6,16,2,1,
/* out0429_em-eta9-phi21*/	7,6,1,11,21,2,1,22,0,2,8,1,8,8,2,5,9,0,1,15,0,3,
/* out0430_em-eta10-phi21*/	9,4,5,6,5,5,9,6,0,3,6,1,2,21,0,1,21,2,2,7,2,1,8,0,8,8,1,6,
/* out0431_em-eta11-phi21*/	9,4,2,2,4,4,1,4,5,10,5,0,14,5,1,2,5,4,7,5,5,3,7,1,3,7,2,9,
/* out0432_em-eta12-phi21*/	7,4,0,2,4,1,15,4,2,7,5,0,2,5,1,5,7,0,9,7,1,1,
/* out0433_em-eta13-phi21*/	7,3,2,6,3,4,5,3,5,13,4,0,1,1,1,1,6,2,6,7,0,2,
/* out0434_em-eta14-phi21*/	6,2,2,8,3,0,2,3,3,1,3,4,11,6,0,3,6,2,4,
/* out0435_em-eta15-phi21*/	6,2,0,8,2,1,3,2,2,5,2,3,3,0,1,2,6,0,4,
/* out0436_em-eta16-phi21*/	4,1,2,10,2,0,5,0,1,3,5,0,4,
/* out0437_em-eta17-phi21*/	7,1,2,4,1,3,7,1,4,2,0,0,1,0,1,1,5,0,5,5,1,1,
/* out0438_em-eta18-phi21*/	4,0,2,1,0,3,5,1,3,3,1,4,1,
/* out0439_em-eta19-phi21*/	2,0,0,3,0,3,5,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	6,10,0,1,10,1,14,10,2,4,25,2,5,26,0,4,26,2,12,
/* out0444_em-eta4-phi22*/	6,9,1,11,9,2,7,10,0,4,10,1,2,25,0,7,25,2,4,
/* out0445_em-eta5-phi22*/	6,8,1,4,8,2,6,9,0,8,9,1,5,24,0,3,24,2,4,
/* out0446_em-eta6-phi22*/	4,8,0,10,8,1,10,8,2,3,10,0,2,
/* out0447_em-eta7-phi22*/	7,7,0,2,7,1,6,7,2,12,4,1,4,9,2,7,10,0,6,10,2,15,
/* out0448_em-eta8-phi22*/	8,6,2,4,7,0,11,7,1,1,3,1,1,4,1,1,9,0,10,9,1,1,9,2,8,
/* out0449_em-eta9-phi22*/	6,6,0,4,6,1,1,6,2,9,3,1,7,8,2,9,9,0,3,
/* out0450_em-eta10-phi22*/	8,5,2,8,5,5,2,6,0,8,2,1,5,2,2,1,3,0,3,8,0,8,8,2,2,
/* out0451_em-eta11-phi22*/	9,4,2,2,4,3,1,5,2,8,5,3,13,5,4,9,5,5,2,2,0,3,2,1,8,7,2,5,
/* out0452_em-eta12-phi22*/	8,4,0,10,4,2,5,4,3,13,1,1,4,1,2,4,2,0,1,7,0,3,7,2,1,
/* out0453_em-eta13-phi22*/	5,3,2,10,3,3,1,4,0,3,1,0,1,1,1,8,
/* out0454_em-eta14-phi22*/	8,2,3,5,3,3,14,0,1,1,0,2,2,1,0,3,1,1,2,6,0,1,6,2,1,
/* out0455_em-eta15-phi22*/	4,2,0,3,2,3,8,0,1,4,0,2,2,
/* out0456_em-eta16-phi22*/	3,0,0,1,0,1,4,0,2,1,
/* out0457_em-eta17-phi22*/	4,1,2,1,1,3,2,0,0,4,0,1,1,
/* out0458_em-eta18-phi22*/	2,0,3,3,1,3,4,
/* out0459_em-eta19-phi22*/	1,0,3,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	2,10,0,6,10,2,12,
/* out0464_em-eta4-phi23*/	3,9,0,1,9,2,9,10,0,5,
/* out0465_em-eta5-phi23*/	2,8,2,3,9,0,7,
/* out0466_em-eta6-phi23*/	2,8,0,6,8,2,4,
/* out0467_em-eta7-phi23*/	6,7,0,1,7,2,4,4,0,7,4,1,9,4,2,16,10,2,1,
/* out0468_em-eta8-phi23*/	5,7,0,2,3,1,2,3,2,12,4,0,9,4,1,2,
/* out0469_em-eta9-phi23*/	5,6,0,1,6,2,2,3,0,9,3,1,6,3,2,4,
/* out0470_em-eta10-phi23*/	3,2,1,1,2,2,13,3,0,4,
/* out0471_em-eta11-phi23*/	4,5,3,3,2,0,9,2,1,2,2,2,2,
/* out0472_em-eta12-phi23*/	3,4,3,2,1,2,8,2,0,3,
/* out0473_em-eta13-phi23*/	3,1,0,6,1,1,1,1,2,4,
/* out0474_em-eta14-phi23*/	2,0,2,2,1,0,6,
/* out0475_em-eta15-phi23*/	1,0,2,7,
/* out0476_em-eta16-phi23*/	2,0,0,4,0,2,2,
/* out0477_em-eta17-phi23*/	1,0,0,5,
/* out0478_em-eta18-phi23*/	1,0,0,1,
/* out0479_em-eta19-phi23*/	0
};