parameter integer matrixH [0:2448] = {
/* num inputs = 170(in0-in169) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 5 */
//* total number of input in adders 944 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	1, 0, 1, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	0, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	1, 3, 1, 
/* out0033_had-eta13-phi1*/	1, 3, 1, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	1, 1, 1, 
/* out0036_had-eta16-phi1*/	1, 1, 1, 
/* out0037_had-eta17-phi1*/	1, 1, 1, 
/* out0038_had-eta18-phi1*/	1, 0, 1, 
/* out0039_had-eta19-phi1*/	1, 0, 2, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	0, 
/* out0045_had-eta5-phi2*/	1, 27, 6, 
/* out0046_had-eta6-phi2*/	2, 26, 4, 27, 1, 
/* out0047_had-eta7-phi2*/	2, 25, 1, 26, 4, 
/* out0048_had-eta8-phi2*/	1, 25, 5, 
/* out0049_had-eta9-phi2*/	2, 24, 1, 25, 2, 
/* out0050_had-eta10-phi2*/	1, 24, 4, 
/* out0051_had-eta11-phi2*/	1, 24, 2, 
/* out0052_had-eta12-phi2*/	1, 3, 3, 
/* out0053_had-eta13-phi2*/	1, 3, 2, 
/* out0054_had-eta14-phi2*/	2, 1, 1, 3, 1, 
/* out0055_had-eta15-phi2*/	1, 1, 2, 
/* out0056_had-eta16-phi2*/	1, 1, 1, 
/* out0057_had-eta17-phi2*/	1, 1, 1, 
/* out0058_had-eta18-phi2*/	1, 0, 2, 
/* out0059_had-eta19-phi2*/	1, 0, 2, 
/* out0060_had-eta0-phi3*/	1, 125, 3, 
/* out0061_had-eta1-phi3*/	2, 124, 1, 125, 5, 
/* out0062_had-eta2-phi3*/	1, 124, 4, 
/* out0063_had-eta3-phi3*/	3, 36, 6, 123, 2, 124, 3, 
/* out0064_had-eta4-phi3*/	4, 27, 1, 35, 4, 36, 1, 123, 4, 
/* out0065_had-eta5-phi3*/	5, 27, 7, 34, 1, 35, 2, 122, 3, 123, 2, 
/* out0066_had-eta6-phi3*/	4, 26, 4, 27, 1, 34, 3, 122, 5, 
/* out0067_had-eta7-phi3*/	3, 25, 1, 26, 4, 33, 2, 
/* out0068_had-eta8-phi3*/	1, 25, 5, 
/* out0069_had-eta9-phi3*/	3, 24, 1, 25, 2, 32, 1, 
/* out0070_had-eta10-phi3*/	1, 24, 4, 
/* out0071_had-eta11-phi3*/	1, 24, 3, 
/* out0072_had-eta12-phi3*/	1, 3, 3, 
/* out0073_had-eta13-phi3*/	1, 3, 2, 
/* out0074_had-eta14-phi3*/	2, 1, 1, 3, 1, 
/* out0075_had-eta15-phi3*/	1, 1, 2, 
/* out0076_had-eta16-phi3*/	1, 1, 1, 
/* out0077_had-eta17-phi3*/	1, 1, 1, 
/* out0078_had-eta18-phi3*/	1, 0, 2, 
/* out0079_had-eta19-phi3*/	1, 0, 2, 
/* out0080_had-eta0-phi4*/	1, 125, 3, 
/* out0081_had-eta1-phi4*/	2, 124, 1, 125, 5, 
/* out0082_had-eta2-phi4*/	1, 124, 4, 
/* out0083_had-eta3-phi4*/	5, 36, 7, 46, 2, 47, 8, 123, 2, 124, 3, 
/* out0084_had-eta4-phi4*/	4, 35, 6, 36, 2, 46, 3, 123, 4, 
/* out0085_had-eta5-phi4*/	5, 34, 4, 35, 4, 45, 2, 122, 3, 123, 2, 
/* out0086_had-eta6-phi4*/	3, 33, 1, 34, 7, 122, 5, 
/* out0087_had-eta7-phi4*/	1, 33, 7, 
/* out0088_had-eta8-phi4*/	2, 32, 2, 33, 3, 
/* out0089_had-eta9-phi4*/	1, 32, 5, 
/* out0090_had-eta10-phi4*/	3, 9, 1, 24, 1, 32, 2, 
/* out0091_had-eta11-phi4*/	1, 9, 3, 
/* out0092_had-eta12-phi4*/	2, 3, 1, 9, 2, 
/* out0093_had-eta13-phi4*/	2, 3, 1, 8, 1, 
/* out0094_had-eta14-phi4*/	1, 8, 2, 
/* out0095_had-eta15-phi4*/	2, 1, 1, 8, 1, 
/* out0096_had-eta16-phi4*/	1, 1, 1, 
/* out0097_had-eta17-phi4*/	1, 1, 1, 
/* out0098_had-eta18-phi4*/	1, 0, 1, 
/* out0099_had-eta19-phi4*/	1, 0, 2, 
/* out0100_had-eta0-phi5*/	1, 129, 3, 
/* out0101_had-eta1-phi5*/	2, 128, 1, 129, 5, 
/* out0102_had-eta2-phi5*/	2, 58, 1, 128, 4, 
/* out0103_had-eta3-phi5*/	5, 46, 4, 47, 8, 58, 6, 127, 2, 128, 3, 
/* out0104_had-eta4-phi5*/	4, 45, 3, 46, 7, 57, 2, 127, 4, 
/* out0105_had-eta5-phi5*/	3, 45, 10, 126, 3, 127, 2, 
/* out0106_had-eta6-phi5*/	3, 34, 1, 44, 8, 126, 5, 
/* out0107_had-eta7-phi5*/	3, 33, 2, 43, 2, 44, 3, 
/* out0108_had-eta8-phi5*/	3, 32, 1, 33, 1, 43, 4, 
/* out0109_had-eta9-phi5*/	1, 32, 4, 
/* out0110_had-eta10-phi5*/	3, 9, 2, 32, 1, 42, 1, 
/* out0111_had-eta11-phi5*/	1, 9, 3, 
/* out0112_had-eta12-phi5*/	1, 9, 3, 
/* out0113_had-eta13-phi5*/	1, 8, 2, 
/* out0114_had-eta14-phi5*/	1, 8, 2, 
/* out0115_had-eta15-phi5*/	1, 8, 2, 
/* out0116_had-eta16-phi5*/	1, 2, 1, 
/* out0117_had-eta17-phi5*/	1, 2, 1, 
/* out0118_had-eta18-phi5*/	1, 2, 1, 
/* out0119_had-eta19-phi5*/	2, 0, 1, 2, 1, 
/* out0120_had-eta0-phi6*/	1, 129, 3, 
/* out0121_had-eta1-phi6*/	2, 128, 1, 129, 5, 
/* out0122_had-eta2-phi6*/	2, 58, 1, 128, 4, 
/* out0123_had-eta3-phi6*/	5, 57, 2, 58, 8, 100, 5, 127, 2, 128, 3, 
/* out0124_had-eta4-phi6*/	2, 57, 12, 127, 4, 
/* out0125_had-eta5-phi6*/	4, 45, 1, 56, 8, 126, 3, 127, 2, 
/* out0126_had-eta6-phi6*/	4, 44, 4, 55, 2, 56, 2, 126, 5, 
/* out0127_had-eta7-phi6*/	3, 43, 3, 44, 1, 55, 2, 
/* out0128_had-eta8-phi6*/	1, 43, 5, 
/* out0129_had-eta9-phi6*/	2, 42, 4, 43, 1, 
/* out0130_had-eta10-phi6*/	1, 42, 4, 
/* out0131_had-eta11-phi6*/	3, 9, 1, 10, 1, 42, 1, 
/* out0132_had-eta12-phi6*/	2, 9, 1, 10, 2, 
/* out0133_had-eta13-phi6*/	1, 8, 2, 
/* out0134_had-eta14-phi6*/	1, 8, 2, 
/* out0135_had-eta15-phi6*/	1, 8, 1, 
/* out0136_had-eta16-phi6*/	1, 2, 1, 
/* out0137_had-eta17-phi6*/	1, 2, 1, 
/* out0138_had-eta18-phi6*/	1, 2, 1, 
/* out0139_had-eta19-phi6*/	1, 2, 1, 
/* out0140_had-eta0-phi7*/	1, 133, 3, 
/* out0141_had-eta1-phi7*/	2, 132, 1, 133, 5, 
/* out0142_had-eta2-phi7*/	2, 102, 7, 132, 4, 
/* out0143_had-eta3-phi7*/	5, 100, 10, 101, 3, 102, 4, 131, 2, 132, 3, 
/* out0144_had-eta4-phi7*/	3, 99, 10, 100, 1, 131, 4, 
/* out0145_had-eta5-phi7*/	5, 56, 5, 98, 3, 99, 2, 130, 3, 131, 2, 
/* out0146_had-eta6-phi7*/	4, 55, 5, 56, 1, 98, 2, 130, 5, 
/* out0147_had-eta7-phi7*/	2, 54, 1, 55, 5, 
/* out0148_had-eta8-phi7*/	2, 43, 1, 54, 5, 
/* out0149_had-eta9-phi7*/	2, 42, 3, 54, 2, 
/* out0150_had-eta10-phi7*/	1, 42, 3, 
/* out0151_had-eta11-phi7*/	1, 10, 3, 
/* out0152_had-eta12-phi7*/	1, 10, 3, 
/* out0153_had-eta13-phi7*/	1, 10, 1, 
/* out0154_had-eta14-phi7*/	2, 8, 1, 14, 1, 
/* out0155_had-eta15-phi7*/	1, 14, 1, 
/* out0156_had-eta16-phi7*/	1, 2, 1, 
/* out0157_had-eta17-phi7*/	1, 2, 1, 
/* out0158_had-eta18-phi7*/	1, 2, 1, 
/* out0159_had-eta19-phi7*/	1, 2, 1, 
/* out0160_had-eta0-phi8*/	1, 133, 3, 
/* out0161_had-eta1-phi8*/	2, 132, 1, 133, 5, 
/* out0162_had-eta2-phi8*/	2, 102, 3, 132, 4, 
/* out0163_had-eta3-phi8*/	4, 101, 10, 102, 2, 131, 2, 132, 3, 
/* out0164_had-eta4-phi8*/	4, 99, 3, 101, 3, 110, 6, 131, 4, 
/* out0165_had-eta5-phi8*/	5, 98, 7, 99, 1, 110, 2, 130, 3, 131, 2, 
/* out0166_had-eta6-phi8*/	4, 55, 1, 98, 4, 108, 3, 130, 5, 
/* out0167_had-eta7-phi8*/	3, 54, 1, 55, 1, 108, 5, 
/* out0168_had-eta8-phi8*/	1, 54, 5, 
/* out0169_had-eta9-phi8*/	2, 54, 2, 64, 3, 
/* out0170_had-eta10-phi8*/	1, 64, 4, 
/* out0171_had-eta11-phi8*/	2, 10, 2, 64, 1, 
/* out0172_had-eta12-phi8*/	1, 10, 3, 
/* out0173_had-eta13-phi8*/	2, 10, 1, 14, 1, 
/* out0174_had-eta14-phi8*/	1, 14, 2, 
/* out0175_had-eta15-phi8*/	1, 14, 2, 
/* out0176_had-eta16-phi8*/	2, 2, 1, 14, 1, 
/* out0177_had-eta17-phi8*/	1, 2, 1, 
/* out0178_had-eta18-phi8*/	1, 2, 1, 
/* out0179_had-eta19-phi8*/	1, 2, 1, 
/* out0180_had-eta0-phi9*/	1, 137, 3, 
/* out0181_had-eta1-phi9*/	2, 136, 1, 137, 5, 
/* out0182_had-eta2-phi9*/	2, 114, 3, 136, 4, 
/* out0183_had-eta3-phi9*/	4, 112, 10, 114, 2, 135, 2, 136, 3, 
/* out0184_had-eta4-phi9*/	4, 110, 6, 111, 3, 112, 3, 135, 4, 
/* out0185_had-eta5-phi9*/	5, 109, 7, 110, 2, 111, 1, 134, 3, 135, 2, 
/* out0186_had-eta6-phi9*/	4, 66, 1, 108, 3, 109, 4, 134, 5, 
/* out0187_had-eta7-phi9*/	3, 65, 1, 66, 1, 108, 5, 
/* out0188_had-eta8-phi9*/	1, 65, 5, 
/* out0189_had-eta9-phi9*/	2, 64, 3, 65, 2, 
/* out0190_had-eta10-phi9*/	1, 64, 4, 
/* out0191_had-eta11-phi9*/	2, 15, 2, 64, 1, 
/* out0192_had-eta12-phi9*/	1, 15, 3, 
/* out0193_had-eta13-phi9*/	2, 14, 1, 15, 1, 
/* out0194_had-eta14-phi9*/	1, 14, 2, 
/* out0195_had-eta15-phi9*/	1, 14, 2, 
/* out0196_had-eta16-phi9*/	2, 14, 1, 18, 1, 
/* out0197_had-eta17-phi9*/	1, 18, 1, 
/* out0198_had-eta18-phi9*/	1, 18, 1, 
/* out0199_had-eta19-phi9*/	1, 18, 1, 
/* out0200_had-eta0-phi10*/	1, 137, 3, 
/* out0201_had-eta1-phi10*/	2, 136, 1, 137, 5, 
/* out0202_had-eta2-phi10*/	2, 114, 7, 136, 4, 
/* out0203_had-eta3-phi10*/	5, 112, 3, 113, 10, 114, 4, 135, 2, 136, 3, 
/* out0204_had-eta4-phi10*/	3, 111, 10, 113, 1, 135, 4, 
/* out0205_had-eta5-phi10*/	5, 67, 5, 109, 3, 111, 2, 134, 3, 135, 2, 
/* out0206_had-eta6-phi10*/	4, 66, 5, 67, 1, 109, 2, 134, 5, 
/* out0207_had-eta7-phi10*/	2, 65, 1, 66, 5, 
/* out0208_had-eta8-phi10*/	2, 65, 5, 77, 1, 
/* out0209_had-eta9-phi10*/	2, 65, 2, 76, 3, 
/* out0210_had-eta10-phi10*/	1, 76, 3, 
/* out0211_had-eta11-phi10*/	1, 15, 3, 
/* out0212_had-eta12-phi10*/	1, 15, 3, 
/* out0213_had-eta13-phi10*/	1, 15, 1, 
/* out0214_had-eta14-phi10*/	2, 14, 1, 19, 1, 
/* out0215_had-eta15-phi10*/	1, 14, 1, 
/* out0216_had-eta16-phi10*/	1, 18, 1, 
/* out0217_had-eta17-phi10*/	1, 18, 1, 
/* out0218_had-eta18-phi10*/	1, 18, 1, 
/* out0219_had-eta19-phi10*/	1, 18, 1, 
/* out0220_had-eta0-phi11*/	1, 141, 3, 
/* out0221_had-eta1-phi11*/	2, 140, 1, 141, 5, 
/* out0222_had-eta2-phi11*/	2, 69, 1, 140, 4, 
/* out0223_had-eta3-phi11*/	5, 68, 2, 69, 8, 113, 5, 139, 2, 140, 3, 
/* out0224_had-eta4-phi11*/	2, 68, 12, 139, 4, 
/* out0225_had-eta5-phi11*/	4, 67, 8, 79, 1, 138, 3, 139, 2, 
/* out0226_had-eta6-phi11*/	4, 66, 2, 67, 2, 78, 4, 138, 5, 
/* out0227_had-eta7-phi11*/	3, 66, 2, 77, 3, 78, 1, 
/* out0228_had-eta8-phi11*/	1, 77, 5, 
/* out0229_had-eta9-phi11*/	2, 76, 4, 77, 1, 
/* out0230_had-eta10-phi11*/	1, 76, 4, 
/* out0231_had-eta11-phi11*/	3, 15, 1, 20, 1, 76, 1, 
/* out0232_had-eta12-phi11*/	2, 15, 2, 20, 1, 
/* out0233_had-eta13-phi11*/	1, 19, 2, 
/* out0234_had-eta14-phi11*/	1, 19, 2, 
/* out0235_had-eta15-phi11*/	1, 19, 1, 
/* out0236_had-eta16-phi11*/	1, 18, 1, 
/* out0237_had-eta17-phi11*/	1, 18, 1, 
/* out0238_had-eta18-phi11*/	1, 18, 1, 
/* out0239_had-eta19-phi11*/	1, 18, 1, 
/* out0240_had-eta0-phi12*/	1, 141, 3, 
/* out0241_had-eta1-phi12*/	2, 140, 1, 141, 5, 
/* out0242_had-eta2-phi12*/	2, 69, 1, 140, 4, 
/* out0243_had-eta3-phi12*/	5, 69, 6, 80, 4, 81, 8, 139, 2, 140, 3, 
/* out0244_had-eta4-phi12*/	4, 68, 2, 79, 3, 80, 7, 139, 4, 
/* out0245_had-eta5-phi12*/	3, 79, 10, 138, 3, 139, 2, 
/* out0246_had-eta6-phi12*/	3, 78, 8, 90, 1, 138, 5, 
/* out0247_had-eta7-phi12*/	3, 77, 2, 78, 3, 89, 2, 
/* out0248_had-eta8-phi12*/	3, 77, 4, 88, 1, 89, 1, 
/* out0249_had-eta9-phi12*/	1, 88, 4, 
/* out0250_had-eta10-phi12*/	3, 20, 2, 76, 1, 88, 1, 
/* out0251_had-eta11-phi12*/	1, 20, 3, 
/* out0252_had-eta12-phi12*/	1, 20, 3, 
/* out0253_had-eta13-phi12*/	1, 19, 2, 
/* out0254_had-eta14-phi12*/	1, 19, 2, 
/* out0255_had-eta15-phi12*/	1, 19, 2, 
/* out0256_had-eta16-phi12*/	1, 18, 1, 
/* out0257_had-eta17-phi12*/	1, 18, 1, 
/* out0258_had-eta18-phi12*/	1, 18, 1, 
/* out0259_had-eta19-phi12*/	2, 4, 1, 18, 1, 
/* out0260_had-eta0-phi13*/	1, 145, 3, 
/* out0261_had-eta1-phi13*/	2, 144, 1, 145, 5, 
/* out0262_had-eta2-phi13*/	1, 144, 4, 
/* out0263_had-eta3-phi13*/	5, 80, 2, 81, 8, 92, 7, 143, 2, 144, 3, 
/* out0264_had-eta4-phi13*/	4, 80, 3, 91, 7, 92, 2, 143, 4, 
/* out0265_had-eta5-phi13*/	5, 79, 2, 90, 4, 91, 3, 142, 3, 143, 2, 
/* out0266_had-eta6-phi13*/	3, 89, 1, 90, 7, 142, 5, 
/* out0267_had-eta7-phi13*/	1, 89, 7, 
/* out0268_had-eta8-phi13*/	2, 88, 2, 89, 3, 
/* out0269_had-eta9-phi13*/	1, 88, 5, 
/* out0270_had-eta10-phi13*/	2, 20, 1, 88, 2, 
/* out0271_had-eta11-phi13*/	1, 20, 3, 
/* out0272_had-eta12-phi13*/	2, 7, 1, 20, 2, 
/* out0273_had-eta13-phi13*/	2, 7, 1, 19, 1, 
/* out0274_had-eta14-phi13*/	1, 19, 2, 
/* out0275_had-eta15-phi13*/	2, 6, 1, 19, 1, 
/* out0276_had-eta16-phi13*/	1, 6, 1, 
/* out0277_had-eta17-phi13*/	1, 6, 1, 
/* out0278_had-eta18-phi13*/	1, 4, 1, 
/* out0279_had-eta19-phi13*/	1, 4, 2, 
/* out0280_had-eta0-phi14*/	1, 145, 3, 
/* out0281_had-eta1-phi14*/	2, 144, 1, 145, 5, 
/* out0282_had-eta2-phi14*/	1, 144, 4, 
/* out0283_had-eta3-phi14*/	3, 92, 6, 143, 2, 144, 3, 
/* out0284_had-eta4-phi14*/	3, 91, 4, 92, 1, 143, 4, 
/* out0285_had-eta5-phi14*/	5, 31, 6, 90, 1, 91, 2, 142, 3, 143, 2, 
/* out0286_had-eta6-phi14*/	4, 30, 4, 31, 1, 90, 3, 142, 5, 
/* out0287_had-eta7-phi14*/	3, 29, 1, 30, 4, 89, 2, 
/* out0288_had-eta8-phi14*/	1, 29, 5, 
/* out0289_had-eta9-phi14*/	3, 28, 1, 29, 2, 88, 1, 
/* out0290_had-eta10-phi14*/	1, 28, 4, 
/* out0291_had-eta11-phi14*/	1, 28, 2, 
/* out0292_had-eta12-phi14*/	1, 7, 3, 
/* out0293_had-eta13-phi14*/	1, 7, 2, 
/* out0294_had-eta14-phi14*/	2, 6, 1, 7, 1, 
/* out0295_had-eta15-phi14*/	1, 6, 2, 
/* out0296_had-eta16-phi14*/	1, 6, 1, 
/* out0297_had-eta17-phi14*/	1, 6, 1, 
/* out0298_had-eta18-phi14*/	1, 4, 2, 
/* out0299_had-eta19-phi14*/	1, 4, 2, 
/* out0300_had-eta0-phi15*/	1, 149, 3, 
/* out0301_had-eta1-phi15*/	2, 148, 1, 149, 5, 
/* out0302_had-eta2-phi15*/	1, 148, 4, 
/* out0303_had-eta3-phi15*/	3, 41, 6, 147, 2, 148, 3, 
/* out0304_had-eta4-phi15*/	4, 31, 1, 40, 4, 41, 1, 147, 4, 
/* out0305_had-eta5-phi15*/	5, 31, 7, 39, 1, 40, 2, 146, 3, 147, 2, 
/* out0306_had-eta6-phi15*/	4, 30, 4, 31, 1, 39, 3, 146, 5, 
/* out0307_had-eta7-phi15*/	3, 29, 1, 30, 4, 38, 2, 
/* out0308_had-eta8-phi15*/	1, 29, 5, 
/* out0309_had-eta9-phi15*/	3, 28, 1, 29, 2, 37, 1, 
/* out0310_had-eta10-phi15*/	1, 28, 4, 
/* out0311_had-eta11-phi15*/	1, 28, 3, 
/* out0312_had-eta12-phi15*/	1, 7, 3, 
/* out0313_had-eta13-phi15*/	1, 7, 2, 
/* out0314_had-eta14-phi15*/	2, 6, 1, 7, 1, 
/* out0315_had-eta15-phi15*/	1, 6, 2, 
/* out0316_had-eta16-phi15*/	1, 6, 1, 
/* out0317_had-eta17-phi15*/	1, 6, 1, 
/* out0318_had-eta18-phi15*/	1, 4, 2, 
/* out0319_had-eta19-phi15*/	1, 4, 2, 
/* out0320_had-eta0-phi16*/	1, 149, 3, 
/* out0321_had-eta1-phi16*/	2, 148, 1, 149, 5, 
/* out0322_had-eta2-phi16*/	1, 148, 4, 
/* out0323_had-eta3-phi16*/	5, 41, 7, 52, 2, 53, 8, 147, 2, 148, 3, 
/* out0324_had-eta4-phi16*/	4, 40, 6, 41, 2, 52, 3, 147, 4, 
/* out0325_had-eta5-phi16*/	5, 39, 4, 40, 4, 51, 2, 146, 3, 147, 2, 
/* out0326_had-eta6-phi16*/	3, 38, 1, 39, 7, 146, 5, 
/* out0327_had-eta7-phi16*/	1, 38, 7, 
/* out0328_had-eta8-phi16*/	2, 37, 2, 38, 3, 
/* out0329_had-eta9-phi16*/	1, 37, 5, 
/* out0330_had-eta10-phi16*/	3, 13, 1, 28, 1, 37, 2, 
/* out0331_had-eta11-phi16*/	1, 13, 3, 
/* out0332_had-eta12-phi16*/	2, 7, 1, 13, 2, 
/* out0333_had-eta13-phi16*/	2, 7, 1, 11, 1, 
/* out0334_had-eta14-phi16*/	1, 11, 2, 
/* out0335_had-eta15-phi16*/	2, 6, 1, 11, 1, 
/* out0336_had-eta16-phi16*/	1, 6, 1, 
/* out0337_had-eta17-phi16*/	1, 6, 1, 
/* out0338_had-eta18-phi16*/	1, 4, 1, 
/* out0339_had-eta19-phi16*/	1, 4, 2, 
/* out0340_had-eta0-phi17*/	1, 153, 3, 
/* out0341_had-eta1-phi17*/	2, 152, 1, 153, 5, 
/* out0342_had-eta2-phi17*/	2, 63, 1, 152, 4, 
/* out0343_had-eta3-phi17*/	5, 52, 4, 53, 8, 63, 6, 151, 2, 152, 3, 
/* out0344_had-eta4-phi17*/	4, 51, 3, 52, 7, 62, 2, 151, 4, 
/* out0345_had-eta5-phi17*/	3, 51, 10, 150, 3, 151, 2, 
/* out0346_had-eta6-phi17*/	3, 39, 1, 50, 8, 150, 5, 
/* out0347_had-eta7-phi17*/	3, 38, 2, 49, 2, 50, 3, 
/* out0348_had-eta8-phi17*/	3, 37, 1, 38, 1, 49, 4, 
/* out0349_had-eta9-phi17*/	1, 37, 4, 
/* out0350_had-eta10-phi17*/	3, 13, 2, 37, 1, 48, 1, 
/* out0351_had-eta11-phi17*/	1, 13, 3, 
/* out0352_had-eta12-phi17*/	1, 13, 3, 
/* out0353_had-eta13-phi17*/	1, 11, 2, 
/* out0354_had-eta14-phi17*/	1, 11, 2, 
/* out0355_had-eta15-phi17*/	1, 11, 2, 
/* out0356_had-eta16-phi17*/	1, 5, 1, 
/* out0357_had-eta17-phi17*/	1, 5, 1, 
/* out0358_had-eta18-phi17*/	1, 5, 1, 
/* out0359_had-eta19-phi17*/	2, 4, 1, 5, 1, 
/* out0360_had-eta0-phi18*/	1, 153, 3, 
/* out0361_had-eta1-phi18*/	2, 152, 1, 153, 5, 
/* out0362_had-eta2-phi18*/	2, 63, 1, 152, 4, 
/* out0363_had-eta3-phi18*/	5, 62, 2, 63, 8, 106, 5, 151, 2, 152, 3, 
/* out0364_had-eta4-phi18*/	2, 62, 12, 151, 4, 
/* out0365_had-eta5-phi18*/	4, 51, 1, 61, 8, 150, 3, 151, 2, 
/* out0366_had-eta6-phi18*/	4, 50, 4, 60, 2, 61, 2, 150, 5, 
/* out0367_had-eta7-phi18*/	3, 49, 3, 50, 1, 60, 2, 
/* out0368_had-eta8-phi18*/	1, 49, 5, 
/* out0369_had-eta9-phi18*/	2, 48, 4, 49, 1, 
/* out0370_had-eta10-phi18*/	1, 48, 4, 
/* out0371_had-eta11-phi18*/	3, 12, 1, 13, 1, 48, 1, 
/* out0372_had-eta12-phi18*/	2, 12, 2, 13, 1, 
/* out0373_had-eta13-phi18*/	1, 11, 2, 
/* out0374_had-eta14-phi18*/	1, 11, 2, 
/* out0375_had-eta15-phi18*/	1, 11, 1, 
/* out0376_had-eta16-phi18*/	1, 5, 1, 
/* out0377_had-eta17-phi18*/	1, 5, 1, 
/* out0378_had-eta18-phi18*/	1, 5, 1, 
/* out0379_had-eta19-phi18*/	1, 5, 1, 
/* out0380_had-eta0-phi19*/	1, 157, 3, 
/* out0381_had-eta1-phi19*/	2, 156, 1, 157, 5, 
/* out0382_had-eta2-phi19*/	2, 107, 7, 156, 4, 
/* out0383_had-eta3-phi19*/	5, 105, 3, 106, 10, 107, 4, 155, 2, 156, 3, 
/* out0384_had-eta4-phi19*/	3, 104, 10, 106, 1, 155, 4, 
/* out0385_had-eta5-phi19*/	5, 61, 5, 103, 3, 104, 2, 154, 3, 155, 2, 
/* out0386_had-eta6-phi19*/	4, 60, 5, 61, 1, 103, 2, 154, 5, 
/* out0387_had-eta7-phi19*/	2, 59, 1, 60, 5, 
/* out0388_had-eta8-phi19*/	2, 49, 1, 59, 5, 
/* out0389_had-eta9-phi19*/	2, 48, 3, 59, 2, 
/* out0390_had-eta10-phi19*/	1, 48, 3, 
/* out0391_had-eta11-phi19*/	1, 12, 3, 
/* out0392_had-eta12-phi19*/	1, 12, 3, 
/* out0393_had-eta13-phi19*/	1, 12, 1, 
/* out0394_had-eta14-phi19*/	2, 11, 1, 16, 1, 
/* out0395_had-eta15-phi19*/	1, 16, 1, 
/* out0396_had-eta16-phi19*/	1, 5, 1, 
/* out0397_had-eta17-phi19*/	1, 5, 1, 
/* out0398_had-eta18-phi19*/	1, 5, 1, 
/* out0399_had-eta19-phi19*/	1, 5, 1, 
/* out0400_had-eta0-phi20*/	1, 157, 3, 
/* out0401_had-eta1-phi20*/	2, 156, 1, 157, 5, 
/* out0402_had-eta2-phi20*/	2, 107, 3, 156, 4, 
/* out0403_had-eta3-phi20*/	4, 105, 10, 107, 2, 155, 2, 156, 3, 
/* out0404_had-eta4-phi20*/	4, 104, 3, 105, 3, 119, 6, 155, 4, 
/* out0405_had-eta5-phi20*/	5, 103, 7, 104, 1, 119, 2, 154, 3, 155, 2, 
/* out0406_had-eta6-phi20*/	4, 60, 1, 103, 4, 115, 3, 154, 5, 
/* out0407_had-eta7-phi20*/	3, 59, 1, 60, 1, 115, 5, 
/* out0408_had-eta8-phi20*/	1, 59, 5, 
/* out0409_had-eta9-phi20*/	2, 59, 2, 70, 3, 
/* out0410_had-eta10-phi20*/	1, 70, 4, 
/* out0411_had-eta11-phi20*/	2, 12, 2, 70, 1, 
/* out0412_had-eta12-phi20*/	1, 12, 3, 
/* out0413_had-eta13-phi20*/	2, 12, 1, 16, 1, 
/* out0414_had-eta14-phi20*/	1, 16, 2, 
/* out0415_had-eta15-phi20*/	1, 16, 2, 
/* out0416_had-eta16-phi20*/	2, 5, 1, 16, 1, 
/* out0417_had-eta17-phi20*/	1, 5, 1, 
/* out0418_had-eta18-phi20*/	1, 5, 1, 
/* out0419_had-eta19-phi20*/	1, 5, 1, 
/* out0420_had-eta0-phi21*/	1, 161, 3, 
/* out0421_had-eta1-phi21*/	2, 160, 1, 161, 5, 
/* out0422_had-eta2-phi21*/	2, 121, 3, 160, 4, 
/* out0423_had-eta3-phi21*/	4, 120, 10, 121, 2, 159, 2, 160, 3, 
/* out0424_had-eta4-phi21*/	4, 117, 3, 119, 6, 120, 3, 159, 4, 
/* out0425_had-eta5-phi21*/	5, 116, 7, 117, 1, 119, 2, 158, 3, 159, 2, 
/* out0426_had-eta6-phi21*/	4, 72, 1, 115, 3, 116, 4, 158, 5, 
/* out0427_had-eta7-phi21*/	3, 71, 1, 72, 1, 115, 5, 
/* out0428_had-eta8-phi21*/	1, 71, 5, 
/* out0429_had-eta9-phi21*/	2, 70, 3, 71, 2, 
/* out0430_had-eta10-phi21*/	1, 70, 4, 
/* out0431_had-eta11-phi21*/	2, 17, 2, 70, 1, 
/* out0432_had-eta12-phi21*/	1, 17, 3, 
/* out0433_had-eta13-phi21*/	2, 16, 1, 17, 1, 
/* out0434_had-eta14-phi21*/	1, 16, 2, 
/* out0435_had-eta15-phi21*/	1, 16, 2, 
/* out0436_had-eta16-phi21*/	2, 16, 1, 21, 1, 
/* out0437_had-eta17-phi21*/	1, 21, 1, 
/* out0438_had-eta18-phi21*/	1, 21, 1, 
/* out0439_had-eta19-phi21*/	1, 21, 1, 
/* out0440_had-eta0-phi22*/	1, 161, 3, 
/* out0441_had-eta1-phi22*/	2, 160, 1, 161, 5, 
/* out0442_had-eta2-phi22*/	2, 121, 7, 160, 4, 
/* out0443_had-eta3-phi22*/	5, 118, 10, 120, 3, 121, 4, 159, 2, 160, 3, 
/* out0444_had-eta4-phi22*/	3, 117, 10, 118, 1, 159, 4, 
/* out0445_had-eta5-phi22*/	5, 73, 5, 116, 3, 117, 2, 158, 3, 159, 2, 
/* out0446_had-eta6-phi22*/	4, 72, 5, 73, 1, 116, 2, 158, 5, 
/* out0447_had-eta7-phi22*/	2, 71, 1, 72, 5, 
/* out0448_had-eta8-phi22*/	2, 71, 5, 83, 1, 
/* out0449_had-eta9-phi22*/	2, 71, 2, 82, 3, 
/* out0450_had-eta10-phi22*/	1, 82, 3, 
/* out0451_had-eta11-phi22*/	1, 17, 3, 
/* out0452_had-eta12-phi22*/	1, 17, 3, 
/* out0453_had-eta13-phi22*/	1, 17, 1, 
/* out0454_had-eta14-phi22*/	2, 16, 1, 22, 1, 
/* out0455_had-eta15-phi22*/	1, 16, 1, 
/* out0456_had-eta16-phi22*/	1, 21, 1, 
/* out0457_had-eta17-phi22*/	1, 21, 1, 
/* out0458_had-eta18-phi22*/	1, 21, 1, 
/* out0459_had-eta19-phi22*/	1, 21, 1, 
/* out0460_had-eta0-phi23*/	1, 165, 3, 
/* out0461_had-eta1-phi23*/	2, 164, 1, 165, 5, 
/* out0462_had-eta2-phi23*/	2, 75, 1, 164, 4, 
/* out0463_had-eta3-phi23*/	5, 74, 2, 75, 8, 118, 5, 163, 2, 164, 3, 
/* out0464_had-eta4-phi23*/	2, 74, 12, 163, 4, 
/* out0465_had-eta5-phi23*/	4, 73, 8, 85, 1, 162, 3, 163, 2, 
/* out0466_had-eta6-phi23*/	4, 72, 2, 73, 2, 84, 4, 162, 5, 
/* out0467_had-eta7-phi23*/	3, 72, 2, 83, 3, 84, 1, 
/* out0468_had-eta8-phi23*/	1, 83, 5, 
/* out0469_had-eta9-phi23*/	2, 82, 4, 83, 1, 
/* out0470_had-eta10-phi23*/	1, 82, 4, 
/* out0471_had-eta11-phi23*/	3, 17, 1, 23, 1, 82, 1, 
/* out0472_had-eta12-phi23*/	2, 17, 2, 23, 1, 
/* out0473_had-eta13-phi23*/	1, 22, 2, 
/* out0474_had-eta14-phi23*/	1, 22, 2, 
/* out0475_had-eta15-phi23*/	1, 22, 1, 
/* out0476_had-eta16-phi23*/	1, 21, 1, 
/* out0477_had-eta17-phi23*/	1, 21, 1, 
/* out0478_had-eta18-phi23*/	1, 21, 1, 
/* out0479_had-eta19-phi23*/	1, 21, 1, 
/* out0480_had-eta0-phi24*/	1, 165, 3, 
/* out0481_had-eta1-phi24*/	2, 164, 1, 165, 5, 
/* out0482_had-eta2-phi24*/	2, 75, 1, 164, 4, 
/* out0483_had-eta3-phi24*/	5, 75, 6, 86, 4, 87, 8, 163, 2, 164, 3, 
/* out0484_had-eta4-phi24*/	4, 74, 2, 85, 3, 86, 7, 163, 4, 
/* out0485_had-eta5-phi24*/	3, 85, 10, 162, 3, 163, 2, 
/* out0486_had-eta6-phi24*/	3, 84, 8, 95, 1, 162, 5, 
/* out0487_had-eta7-phi24*/	3, 83, 2, 84, 3, 94, 2, 
/* out0488_had-eta8-phi24*/	3, 83, 4, 93, 1, 94, 1, 
/* out0489_had-eta9-phi24*/	1, 93, 4, 
/* out0490_had-eta10-phi24*/	3, 23, 2, 82, 1, 93, 1, 
/* out0491_had-eta11-phi24*/	1, 23, 3, 
/* out0492_had-eta12-phi24*/	1, 23, 3, 
/* out0493_had-eta13-phi24*/	1, 22, 2, 
/* out0494_had-eta14-phi24*/	1, 22, 2, 
/* out0495_had-eta15-phi24*/	1, 22, 2, 
/* out0496_had-eta16-phi24*/	1, 21, 1, 
/* out0497_had-eta17-phi24*/	1, 21, 1, 
/* out0498_had-eta18-phi24*/	1, 21, 1, 
/* out0499_had-eta19-phi24*/	1, 21, 1, 
/* out0500_had-eta0-phi25*/	1, 169, 3, 
/* out0501_had-eta1-phi25*/	2, 168, 1, 169, 5, 
/* out0502_had-eta2-phi25*/	1, 168, 4, 
/* out0503_had-eta3-phi25*/	5, 86, 2, 87, 8, 97, 7, 167, 2, 168, 3, 
/* out0504_had-eta4-phi25*/	4, 86, 3, 96, 6, 97, 2, 167, 4, 
/* out0505_had-eta5-phi25*/	5, 85, 2, 95, 4, 96, 4, 166, 3, 167, 2, 
/* out0506_had-eta6-phi25*/	3, 94, 1, 95, 7, 166, 5, 
/* out0507_had-eta7-phi25*/	1, 94, 7, 
/* out0508_had-eta8-phi25*/	2, 93, 2, 94, 3, 
/* out0509_had-eta9-phi25*/	1, 93, 5, 
/* out0510_had-eta10-phi25*/	2, 23, 1, 93, 2, 
/* out0511_had-eta11-phi25*/	1, 23, 3, 
/* out0512_had-eta12-phi25*/	1, 23, 2, 
/* out0513_had-eta13-phi25*/	1, 22, 1, 
/* out0514_had-eta14-phi25*/	1, 22, 2, 
/* out0515_had-eta15-phi25*/	1, 22, 1, 
/* out0516_had-eta16-phi25*/	0, 
/* out0517_had-eta17-phi25*/	0, 
/* out0518_had-eta18-phi25*/	0, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	1, 169, 3, 
/* out0521_had-eta1-phi26*/	2, 168, 1, 169, 5, 
/* out0522_had-eta2-phi26*/	1, 168, 4, 
/* out0523_had-eta3-phi26*/	3, 97, 6, 167, 2, 168, 3, 
/* out0524_had-eta4-phi26*/	3, 96, 4, 97, 1, 167, 4, 
/* out0525_had-eta5-phi26*/	4, 95, 1, 96, 2, 166, 3, 167, 2, 
/* out0526_had-eta6-phi26*/	2, 95, 3, 166, 5, 
/* out0527_had-eta7-phi26*/	1, 94, 2, 
/* out0528_had-eta8-phi26*/	0, 
/* out0529_had-eta9-phi26*/	1, 93, 1, 
/* out0530_had-eta10-phi26*/	0, 
/* out0531_had-eta11-phi26*/	0, 
/* out0532_had-eta12-phi26*/	0, 
/* out0533_had-eta13-phi26*/	0, 
/* out0534_had-eta14-phi26*/	0, 
/* out0535_had-eta15-phi26*/	0, 
/* out0536_had-eta16-phi26*/	0, 
/* out0537_had-eta17-phi26*/	0, 
/* out0538_had-eta18-phi26*/	0, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	0, 
/* out0550_had-eta10-phi27*/	0, 
/* out0551_had-eta11-phi27*/	0, 
/* out0552_had-eta12-phi27*/	0, 
/* out0553_had-eta13-phi27*/	0, 
/* out0554_had-eta14-phi27*/	0, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	0, 
/* out0557_had-eta17-phi27*/	0, 
/* out0558_had-eta18-phi27*/	0, 
/* out0559_had-eta19-phi27*/	0, 
};