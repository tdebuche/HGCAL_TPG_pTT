parameter integer matrixH [0:8180] = {
/* num inputs = 302(in0-in301) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 11 */
//* total number of input in adders 2566 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	1,142,0,16,
/* out0002_em-eta2-phi0*/	2,141,0,1,142,1,16,
/* out0003_em-eta3-phi0*/	7,134,1,4,136,0,1,136,1,8,137,0,15,137,2,9,141,0,15,141,1,3,
/* out0004_em-eta4-phi0*/	9,133,1,6,133,2,3,134,0,2,134,1,5,136,0,15,136,1,8,136,2,16,140,0,3,141,1,13,
/* out0005_em-eta5-phi0*/	7,132,1,15,132,2,2,133,0,11,133,1,10,133,2,3,140,0,13,140,1,5,
/* out0006_em-eta6-phi0*/	7,94,0,3,132,0,11,132,1,1,132,2,14,133,0,1,139,0,6,140,1,11,
/* out0007_em-eta7-phi0*/	5,93,1,12,93,2,2,132,0,5,139,0,10,139,1,7,
/* out0008_em-eta8-phi0*/	6,92,1,15,92,2,2,93,0,8,93,1,4,139,1,9,139,2,7,
/* out0009_em-eta9-phi0*/	5,92,0,1,92,1,1,92,2,11,138,0,6,139,2,9,
/* out0010_em-eta10-phi0*/	6,34,4,3,35,1,6,92,0,8,92,2,1,138,0,10,138,1,12,
/* out0011_em-eta11-phi0*/	8,34,0,2,34,1,16,34,2,6,35,0,2,35,1,8,92,0,6,127,2,10,138,1,4,
/* out0012_em-eta12-phi0*/	9,32,5,1,33,5,5,34,0,14,34,2,2,34,3,6,126,0,4,126,1,1,127,1,1,127,2,1,
/* out0013_em-eta13-phi0*/	7,32,5,15,33,0,1,33,2,4,33,3,1,33,4,8,33,5,11,126,0,9,
/* out0014_em-eta14-phi0*/	8,32,2,8,32,3,2,33,0,15,33,3,2,33,4,8,125,0,1,126,0,1,126,2,1,
/* out0015_em-eta15-phi0*/	6,32,0,8,32,1,16,32,2,8,32,3,7,42,4,1,125,0,6,
/* out0016_em-eta16-phi0*/	3,32,0,8,42,4,12,125,0,4,
/* out0017_em-eta17-phi0*/	3,42,4,2,43,1,9,124,0,1,
/* out0018_em-eta18-phi0*/	3,42,1,4,43,1,5,124,0,4,
/* out0019_em-eta19-phi0*/	1,42,1,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	1,142,3,16,
/* out0022_em-eta2-phi1*/	6,135,1,3,135,2,7,137,0,1,137,2,1,141,3,1,142,2,16,
/* out0023_em-eta3-phi1*/	9,96,0,1,134,1,5,134,2,10,135,0,12,135,1,13,135,2,2,137,2,6,141,2,3,141,3,15,
/* out0024_em-eta4-phi1*/	8,95,0,1,95,1,5,133,2,3,134,0,14,134,1,2,134,2,6,140,3,3,141,2,13,
/* out0025_em-eta5-phi1*/	6,94,1,6,95,0,10,133,0,4,133,2,7,140,2,5,140,3,13,
/* out0026_em-eta6-phi1*/	5,94,0,10,94,1,8,94,2,4,139,5,6,140,2,11,
/* out0027_em-eta7-phi1*/	6,93,2,11,94,0,3,94,2,2,104,0,1,139,4,7,139,5,10,
/* out0028_em-eta8-phi1*/	5,93,0,8,93,2,3,103,1,3,139,3,7,139,4,9,
/* out0029_em-eta9-phi1*/	5,92,2,1,103,0,1,103,1,11,138,3,6,139,3,9,
/* out0030_em-eta10-phi1*/	9,34,4,13,34,5,8,35,1,1,92,0,1,92,2,1,103,0,3,103,1,1,138,2,12,138,3,10,
/* out0031_em-eta11-phi1*/	9,34,2,4,34,5,3,35,0,14,35,1,1,35,4,11,35,5,1,127,1,11,127,2,5,138,2,4,
/* out0032_em-eta12-phi1*/	7,34,2,4,34,3,8,35,3,12,35,4,5,122,0,1,126,1,10,127,1,3,
/* out0033_em-eta13-phi1*/	8,33,2,11,34,3,2,35,3,1,44,1,6,45,1,3,126,0,2,126,1,2,126,2,6,
/* out0034_em-eta14-phi1*/	7,32,3,1,33,2,1,33,3,13,44,0,4,44,1,1,125,1,5,126,2,4,
/* out0035_em-eta15-phi1*/	6,32,3,6,42,5,9,43,5,2,125,0,3,125,1,4,125,2,1,
/* out0036_em-eta16-phi1*/	5,42,4,1,42,5,7,43,0,6,125,0,2,125,2,4,
/* out0037_em-eta17-phi1*/	6,42,2,2,43,0,8,43,1,2,124,0,1,124,1,4,125,2,1,
/* out0038_em-eta18-phi1*/	3,42,1,8,42,2,2,124,0,6,
/* out0039_em-eta19-phi1*/	2,42,0,2,42,1,2,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	1,147,0,16,
/* out0042_em-eta2-phi2*/	5,97,1,4,97,2,5,135,2,4,146,0,1,147,1,16,
/* out0043_em-eta3-phi2*/	9,96,0,4,96,1,16,96,2,4,97,1,1,97,2,10,135,0,4,135,2,3,146,0,15,146,1,3,
/* out0044_em-eta4-phi2*/	7,95,1,10,95,2,3,96,0,11,96,2,5,106,1,3,145,0,3,146,1,13,
/* out0045_em-eta5-phi2*/	7,94,1,1,95,0,5,95,1,1,95,2,13,105,1,6,145,0,13,145,1,5,
/* out0046_em-eta6-phi2*/	7,94,1,1,94,2,9,104,1,2,105,0,3,105,1,8,144,0,6,145,1,11,
/* out0047_em-eta7-phi2*/	6,94,2,1,104,0,6,104,1,11,104,2,1,144,0,10,144,1,7,
/* out0048_em-eta8-phi2*/	5,103,2,6,104,0,9,104,2,1,144,1,9,144,2,7,
/* out0049_em-eta9-phi2*/	5,103,0,4,103,1,1,103,2,7,143,0,6,144,2,9,
/* out0050_em-eta10-phi2*/	6,34,5,4,35,5,1,46,4,10,103,0,7,143,0,10,143,1,12,
/* out0051_em-eta11-phi2*/	9,34,5,1,35,2,6,35,5,14,46,4,5,47,1,8,122,0,7,122,1,7,127,1,1,143,1,4,
/* out0052_em-eta12-phi2*/	9,35,2,10,35,3,3,44,4,10,45,1,4,46,1,1,47,1,1,122,0,8,122,2,3,126,1,2,
/* out0053_em-eta13-phi2*/	8,44,1,5,44,2,5,45,0,6,45,1,9,121,0,5,121,1,1,126,1,1,126,2,4,
/* out0054_em-eta14-phi2*/	7,44,0,8,44,1,4,44,2,5,44,3,3,121,0,5,125,1,3,126,2,1,
/* out0055_em-eta15-phi2*/	6,43,2,1,43,5,10,44,0,4,44,3,2,125,1,4,125,2,3,
/* out0056_em-eta16-phi2*/	4,43,0,1,43,4,9,43,5,4,125,2,6,
/* out0057_em-eta17-phi2*/	4,42,2,7,43,0,1,43,4,4,124,1,6,
/* out0058_em-eta18-phi2*/	6,42,0,3,42,1,1,42,2,4,42,3,2,124,0,3,124,1,2,
/* out0059_em-eta19-phi2*/	1,42,0,7,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	1,147,3,16,
/* out0062_em-eta2-phi3*/	3,97,1,3,146,3,1,147,2,16,
/* out0063_em-eta3-phi3*/	8,96,2,4,97,1,8,97,2,1,107,0,6,107,1,16,107,2,7,146,2,3,146,3,15,
/* out0064_em-eta4-phi3*/	7,96,2,3,106,0,3,106,1,11,106,2,12,107,0,4,145,3,3,146,2,13,
/* out0065_em-eta5-phi3*/	7,105,1,1,105,2,11,106,0,11,106,1,2,115,1,2,145,2,5,145,3,13,
/* out0066_em-eta6-phi3*/	6,105,0,13,105,1,1,105,2,4,114,1,3,144,5,6,145,2,11,
/* out0067_em-eta7-phi3*/	5,104,1,3,104,2,9,114,1,6,144,4,7,144,5,10,
/* out0068_em-eta8-phi3*/	5,104,2,5,113,0,2,113,1,8,144,3,7,144,4,9,
/* out0069_em-eta9-phi3*/	7,46,5,1,47,5,1,103,0,1,103,2,3,113,0,9,143,3,6,144,3,9,
/* out0070_em-eta10-phi3*/	7,46,4,1,46,5,15,47,0,7,47,4,6,47,5,11,143,2,12,143,3,10,
/* out0071_em-eta11-phi3*/	8,46,1,7,46,2,9,47,0,9,47,1,7,47,4,1,122,1,9,122,2,3,143,2,4,
/* out0072_em-eta12-phi3*/	7,44,4,6,44,5,12,46,0,4,46,1,8,121,1,2,122,2,10,123,1,1,
/* out0073_em-eta13-phi3*/	7,44,2,1,44,5,2,45,0,10,45,4,9,45,5,1,121,0,1,121,1,9,
/* out0074_em-eta14-phi3*/	6,44,2,5,44,3,4,45,3,5,45,4,6,121,0,4,121,2,5,
/* out0075_em-eta15-phi3*/	8,43,2,6,44,3,7,45,3,3,120,0,2,120,1,3,121,0,1,121,2,2,125,2,1,
/* out0076_em-eta16-phi3*/	4,43,2,8,43,3,5,43,4,1,120,0,6,
/* out0077_em-eta17-phi3*/	6,42,2,1,42,3,3,43,3,6,43,4,2,120,0,4,124,1,2,
/* out0078_em-eta18-phi3*/	4,42,0,2,42,3,8,124,0,1,124,1,2,
/* out0079_em-eta19-phi3*/	2,0,0,2,42,0,2,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	1,152,0,16,
/* out0082_em-eta2-phi4*/	2,151,0,1,152,1,16,
/* out0083_em-eta3-phi4*/	8,107,0,5,107,2,9,116,1,2,116,2,4,117,1,4,117,2,14,151,0,15,151,1,3,
/* out0084_em-eta4-phi4*/	9,106,0,1,106,2,4,107,0,1,115,2,1,116,0,8,116,1,14,116,2,3,150,0,3,151,1,13,
/* out0085_em-eta5-phi4*/	6,106,0,1,115,0,4,115,1,13,115,2,8,150,0,13,150,1,5,
/* out0086_em-eta6-phi4*/	7,105,2,1,114,1,3,114,2,10,115,0,7,115,1,1,149,0,6,150,1,11,
/* out0087_em-eta7-phi4*/	5,114,0,12,114,1,4,114,2,2,149,0,10,149,1,7,
/* out0088_em-eta8-phi4*/	5,113,1,8,113,2,6,114,0,1,149,1,9,149,2,7,
/* out0089_em-eta9-phi4*/	4,113,0,5,113,2,7,148,0,6,149,2,9,
/* out0090_em-eta10-phi4*/	7,47,2,16,47,3,9,47,4,5,47,5,4,48,0,1,148,0,10,148,1,12,
/* out0091_em-eta11-phi4*/	8,46,0,3,46,2,7,46,3,14,47,3,5,47,4,4,123,1,2,123,2,7,148,1,4,
/* out0092_em-eta12-phi4*/	8,6,5,6,7,5,7,44,5,2,45,5,4,46,0,9,123,0,1,123,1,11,123,2,1,
/* out0093_em-eta13-phi4*/	10,6,4,2,6,5,3,45,2,7,45,4,1,45,5,11,116,0,1,121,1,4,121,2,3,123,0,1,123,1,2,
/* out0094_em-eta14-phi4*/	6,3,2,3,3,5,1,45,2,9,45,3,6,116,0,2,121,2,6,
/* out0095_em-eta15-phi4*/	4,2,5,4,3,5,11,45,3,2,120,1,7,
/* out0096_em-eta16-phi4*/	7,2,4,2,2,5,9,43,2,1,43,3,1,120,0,2,120,1,2,120,2,2,
/* out0097_em-eta17-phi4*/	6,1,1,1,2,4,5,42,3,1,43,3,4,120,0,2,120,2,4,
/* out0098_em-eta18-phi4*/	3,0,0,2,0,1,10,42,3,2,
/* out0099_em-eta19-phi4*/	1,0,0,6,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	1,152,3,16,
/* out0102_em-eta2-phi5*/	2,151,3,1,152,2,16,
/* out0103_em-eta3-phi5*/	5,116,2,3,117,1,12,117,2,2,151,2,3,151,3,15,
/* out0104_em-eta4-phi5*/	6,51,0,8,51,1,4,116,0,8,116,2,6,150,3,3,151,2,13,
/* out0105_em-eta5-phi5*/	8,50,0,1,50,1,2,51,0,8,51,2,4,115,0,3,115,2,7,150,2,5,150,3,13,
/* out0106_em-eta6-phi5*/	7,50,0,14,50,1,1,50,2,2,114,2,2,115,0,2,149,5,6,150,2,11,
/* out0107_em-eta7-phi5*/	8,49,0,6,49,1,4,50,0,1,50,2,2,114,0,3,114,2,2,149,4,7,149,5,10,
/* out0108_em-eta8-phi5*/	5,49,0,10,49,2,3,113,2,1,149,3,7,149,4,9,
/* out0109_em-eta9-phi5*/	6,48,0,6,48,1,4,49,2,1,113,2,2,148,3,6,149,3,9,
/* out0110_em-eta10-phi5*/	4,48,0,8,48,2,2,148,2,12,148,3,10,
/* out0111_em-eta11-phi5*/	10,7,2,16,7,3,4,7,5,1,46,3,2,47,3,2,48,0,1,48,2,2,123,0,1,123,2,7,148,2,4,
/* out0112_em-eta12-phi5*/	6,6,5,3,7,0,7,7,4,11,7,5,8,123,0,11,123,2,1,
/* out0113_em-eta13-phi5*/	7,6,4,11,6,5,4,7,0,5,7,1,3,116,0,1,116,1,7,123,0,2,
/* out0114_em-eta14-phi5*/	5,3,2,13,3,3,4,3,5,1,6,4,3,116,0,9,
/* out0115_em-eta15-phi5*/	5,3,0,2,3,4,11,3,5,3,116,0,3,120,1,3,
/* out0116_em-eta16-phi5*/	6,2,4,1,2,5,3,3,0,9,3,1,1,120,1,1,120,2,6,
/* out0117_em-eta17-phi5*/	4,1,1,2,2,4,8,3,1,3,120,2,4,
/* out0118_em-eta18-phi5*/	4,0,1,5,0,2,7,1,0,4,1,1,9,
/* out0119_em-eta19-phi5*/	4,0,0,6,0,1,1,0,2,5,0,3,2,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	1,157,0,16,
/* out0122_em-eta2-phi6*/	2,156,0,1,157,1,16,
/* out0123_em-eta3-phi6*/	5,59,1,3,60,1,2,60,2,12,156,0,15,156,1,3,
/* out0124_em-eta4-phi6*/	5,51,1,12,59,0,8,59,1,6,155,0,3,156,1,13,
/* out0125_em-eta5-phi6*/	6,50,1,4,51,2,12,58,0,9,58,1,1,155,0,13,155,1,5,
/* out0126_em-eta6-phi6*/	6,50,1,9,50,2,9,57,1,2,58,0,2,154,0,6,155,1,11,
/* out0127_em-eta7-phi6*/	6,49,1,10,50,2,3,57,0,3,57,1,2,154,0,10,154,1,7,
/* out0128_em-eta8-phi6*/	5,49,1,2,49,2,11,56,0,1,154,1,9,154,2,7,
/* out0129_em-eta9-phi6*/	5,48,1,10,49,2,1,56,0,2,153,0,6,154,2,9,
/* out0130_em-eta10-phi6*/	4,48,1,2,48,2,9,153,0,10,153,1,12,
/* out0131_em-eta11-phi6*/	9,6,3,8,7,3,12,7,4,1,18,5,2,19,5,2,48,2,2,118,0,1,118,1,7,153,1,4,
/* out0132_em-eta12-phi6*/	8,6,0,1,6,1,2,6,2,14,6,3,6,7,0,1,7,4,4,118,0,11,118,1,1,
/* out0133_em-eta13-phi6*/	7,6,1,9,6,2,2,7,0,3,7,1,10,116,1,8,116,2,1,118,0,2,
/* out0134_em-eta14-phi6*/	6,2,3,4,3,3,12,3,4,1,7,1,3,116,1,1,116,2,8,
/* out0135_em-eta15-phi6*/	5,2,2,10,2,3,3,3,4,4,115,2,3,116,2,3,
/* out0136_em-eta16-phi6*/	6,2,1,3,2,2,6,3,0,5,3,1,1,115,1,6,115,2,1,
/* out0137_em-eta17-phi6*/	4,0,4,2,2,1,1,3,1,10,115,1,4,
/* out0138_em-eta18-phi6*/	4,0,4,6,0,5,1,1,0,6,1,1,4,
/* out0139_em-eta19-phi6*/	5,0,2,4,0,3,8,1,0,5,1,3,4,1,5,4,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	1,157,3,16,
/* out0142_em-eta2-phi7*/	2,156,3,1,157,2,16,
/* out0143_em-eta3-phi7*/	8,59,1,4,59,2,2,60,1,14,60,2,4,70,0,5,70,1,9,156,2,3,156,3,15,
/* out0144_em-eta4-phi7*/	8,58,1,1,59,0,8,59,1,3,59,2,14,69,0,5,70,0,1,155,3,3,156,2,13,
/* out0145_em-eta5-phi7*/	6,58,0,4,58,1,14,58,2,7,69,0,1,155,2,5,155,3,13,
/* out0146_em-eta6-phi7*/	7,57,1,10,57,2,3,58,0,1,58,2,8,68,1,1,154,5,6,155,2,11,
/* out0147_em-eta7-phi7*/	5,57,0,12,57,1,2,57,2,4,154,4,7,154,5,10,
/* out0148_em-eta8-phi7*/	5,56,0,6,56,1,8,57,0,1,154,3,7,154,4,9,
/* out0149_em-eta9-phi7*/	4,56,0,7,56,2,5,153,3,6,154,3,9,
/* out0150_em-eta10-phi7*/	7,19,2,16,19,3,4,19,4,5,19,5,9,48,2,1,153,2,12,153,3,10,
/* out0151_em-eta11-phi7*/	9,6,3,1,18,4,3,18,5,14,19,0,7,19,4,4,19,5,5,118,1,7,118,2,2,153,2,4,
/* out0152_em-eta12-phi7*/	7,6,0,13,6,3,1,17,2,6,18,4,9,118,0,1,118,1,1,118,2,11,
/* out0153_em-eta13-phi7*/	9,6,0,2,6,1,5,17,2,4,17,5,14,116,2,1,117,1,3,117,2,4,118,0,1,118,2,2,
/* out0154_em-eta14-phi7*/	6,2,3,5,16,4,1,16,5,13,17,5,1,116,2,3,117,1,6,
/* out0155_em-eta15-phi7*/	4,2,0,11,2,3,4,16,4,2,115,2,7,
/* out0156_em-eta16-phi7*/	7,2,0,4,2,1,8,5,2,1,5,5,1,115,0,2,115,1,2,115,2,2,
/* out0157_em-eta17-phi7*/	7,0,4,1,2,1,4,3,1,1,4,5,1,5,5,4,115,0,2,115,1,4,
/* out0158_em-eta18-phi7*/	3,0,4,7,0,5,5,4,5,2,
/* out0159_em-eta19-phi7*/	5,0,3,5,0,5,5,1,0,1,1,3,10,1,5,10,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	1,162,0,16,
/* out0162_em-eta2-phi8*/	3,80,2,3,161,0,1,162,1,16,
/* out0163_em-eta3-phi8*/	7,70,0,6,70,1,7,70,2,16,79,0,4,80,0,9,161,0,15,161,1,3,
/* out0164_em-eta4-phi8*/	7,69,0,6,69,1,15,69,2,5,70,0,4,79,0,3,160,0,3,161,1,13,
/* out0165_em-eta5-phi8*/	7,58,2,1,68,1,11,68,2,1,69,0,4,69,2,9,160,0,13,160,1,5,
/* out0166_em-eta6-phi8*/	7,57,2,3,67,1,1,68,0,13,68,1,4,68,2,1,159,0,6,160,1,11,
/* out0167_em-eta7-phi8*/	5,57,2,6,67,0,2,67,1,10,159,0,10,159,1,7,
/* out0168_em-eta8-phi8*/	5,56,1,8,56,2,2,67,0,5,159,1,9,159,2,7,
/* out0169_em-eta9-phi8*/	7,18,3,1,19,3,1,56,2,9,66,0,1,66,1,3,158,0,6,159,2,9,
/* out0170_em-eta10-phi8*/	7,18,0,1,18,2,7,18,3,15,19,3,11,19,4,6,158,0,10,158,1,12,
/* out0171_em-eta11-phi8*/	8,18,1,7,18,2,9,19,0,9,19,1,7,19,4,1,119,1,3,119,2,9,158,1,4,
/* out0172_em-eta12-phi8*/	7,17,2,5,17,3,12,18,4,4,19,1,8,117,2,2,118,2,1,119,1,10,
/* out0173_em-eta13-phi8*/	8,16,2,3,17,0,2,17,2,1,17,3,2,17,4,16,17,5,1,117,0,1,117,2,9,
/* out0174_em-eta14-phi8*/	6,16,4,3,16,5,3,17,0,11,17,1,3,117,0,4,117,1,5,
/* out0175_em-eta15-phi8*/	9,2,0,1,5,2,6,16,4,10,17,1,1,112,1,1,115,0,2,115,2,3,117,0,1,117,1,2,
/* out0176_em-eta16-phi8*/	4,5,2,8,5,4,1,5,5,5,115,0,6,
/* out0177_em-eta17-phi8*/	6,4,5,3,5,0,1,5,4,2,5,5,6,111,1,2,115,0,4,
/* out0178_em-eta18-phi8*/	4,0,5,1,4,4,2,4,5,8,111,1,3,
/* out0179_em-eta19-phi8*/	5,0,3,1,0,5,4,1,3,2,1,5,2,4,4,2,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	1,162,3,16,
/* out0182_em-eta2-phi9*/	5,80,2,9,120,0,7,120,1,2,161,3,1,162,2,16,
/* out0183_em-eta3-phi9*/	9,79,0,4,79,1,16,79,2,4,80,0,7,80,2,4,120,0,8,120,2,5,161,2,3,161,3,15,
/* out0184_em-eta4-phi9*/	8,69,1,1,69,2,2,78,0,3,78,1,10,79,0,5,79,2,11,160,3,3,161,2,13,
/* out0185_em-eta5-phi9*/	7,68,2,6,77,1,1,78,0,13,78,1,1,78,2,5,160,2,5,160,3,13,
/* out0186_em-eta6-phi9*/	8,67,1,1,67,2,1,68,0,3,68,2,8,77,0,3,77,1,7,159,5,6,160,2,11,
/* out0187_em-eta7-phi9*/	6,67,0,2,67,1,4,67,2,11,77,0,1,159,4,7,159,5,10,
/* out0188_em-eta8-phi9*/	5,66,1,6,67,0,7,67,2,2,159,3,7,159,4,9,
/* out0189_em-eta9-phi9*/	5,66,0,4,66,1,7,66,2,1,158,3,6,159,3,9,
/* out0190_em-eta10-phi9*/	6,18,0,10,20,3,4,21,3,1,66,0,7,158,2,12,158,3,10,
/* out0191_em-eta11-phi9*/	9,18,0,5,18,1,8,20,3,1,21,2,6,21,3,14,114,1,1,119,0,7,119,2,7,158,2,4,
/* out0192_em-eta12-phi9*/	10,16,0,1,16,3,11,17,3,2,18,1,1,19,1,1,21,2,10,21,5,3,113,2,2,119,0,8,119,1,3,
/* out0193_em-eta13-phi9*/	8,16,0,6,16,1,3,16,2,10,16,3,5,113,1,4,113,2,1,117,0,5,117,2,1,
/* out0194_em-eta14-phi9*/	7,16,1,8,16,2,3,17,0,3,17,1,7,112,2,3,113,1,1,117,0,5,
/* out0195_em-eta15-phi9*/	5,5,2,1,5,3,10,17,1,5,112,1,3,112,2,4,
/* out0196_em-eta16-phi9*/	4,4,2,1,5,3,4,5,4,9,112,1,6,
/* out0197_em-eta17-phi9*/	5,4,2,1,5,0,7,5,4,4,111,1,3,111,2,3,
/* out0198_em-eta18-phi9*/	5,4,4,3,4,5,2,5,0,4,5,1,1,111,1,5,
/* out0199_em-eta19-phi9*/	1,4,4,7,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	1,167,0,16,
/* out0202_em-eta2-phi10*/	5,120,1,7,121,0,1,121,2,1,166,0,1,167,1,16,
/* out0203_em-eta3-phi10*/	9,79,2,1,119,1,10,119,2,5,120,0,1,120,1,7,120,2,11,121,0,6,166,0,15,166,1,3,
/* out0204_em-eta4-phi10*/	9,78,1,5,78,2,1,118,0,1,118,1,3,119,0,14,119,1,6,119,2,2,165,0,3,166,1,13,
/* out0205_em-eta5-phi10*/	6,77,1,3,77,2,3,78,2,10,118,0,10,165,0,13,165,1,5,
/* out0206_em-eta6-phi10*/	5,77,0,7,77,1,5,77,2,10,164,0,6,165,1,11,
/* out0207_em-eta7-phi10*/	5,67,2,2,76,1,11,77,0,5,164,0,10,164,1,7,
/* out0208_em-eta8-phi10*/	5,66,2,3,76,0,8,76,1,3,164,1,9,164,2,7,
/* out0209_em-eta9-phi10*/	5,66,0,1,66,2,11,86,1,1,163,0,6,164,2,9,
/* out0210_em-eta10-phi10*/	7,20,0,13,20,1,1,20,3,8,66,0,3,66,2,1,163,0,10,163,1,12,
/* out0211_em-eta11-phi10*/	9,20,1,1,20,2,14,20,3,3,21,0,4,21,3,1,21,4,11,114,0,5,114,1,11,163,1,4,
/* out0212_em-eta12-phi10*/	7,20,5,8,21,0,4,21,4,5,21,5,12,113,2,10,114,1,3,119,0,1,
/* out0213_em-eta13-phi10*/	8,16,0,9,20,5,2,21,5,1,28,5,7,29,5,3,113,0,2,113,1,6,113,2,2,
/* out0214_em-eta14-phi10*/	5,16,1,5,28,4,8,28,5,4,112,2,5,113,1,4,
/* out0215_em-eta15-phi10*/	6,4,3,9,5,3,2,28,4,5,112,0,3,112,1,1,112,2,4,
/* out0216_em-eta16-phi10*/	5,4,0,1,4,2,6,4,3,7,112,0,2,112,1,4,
/* out0217_em-eta17-phi10*/	5,4,1,2,4,2,8,5,0,2,111,2,5,112,1,1,
/* out0218_em-eta18-phi10*/	4,5,0,2,5,1,8,111,1,2,111,2,4,
/* out0219_em-eta19-phi10*/	2,4,4,2,5,1,2,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	1,167,3,16,
/* out0222_em-eta2-phi11*/	2,166,3,1,167,2,16,
/* out0223_em-eta3-phi11*/	7,119,2,4,121,0,9,121,2,15,128,0,1,128,1,7,166,2,3,166,3,15,
/* out0224_em-eta4-phi11*/	7,118,1,9,119,0,2,119,2,5,128,0,15,128,1,1,165,3,3,166,2,13,
/* out0225_em-eta5-phi11*/	6,118,0,5,118,1,4,118,2,16,126,2,2,165,2,5,165,3,13,
/* out0226_em-eta6-phi11*/	5,77,2,3,126,1,3,126,2,14,164,5,6,165,2,11,
/* out0227_em-eta7-phi11*/	5,76,1,2,76,2,12,126,1,4,164,4,7,164,5,10,
/* out0228_em-eta8-phi11*/	5,76,0,8,76,2,4,86,2,2,164,3,7,164,4,9,
/* out0229_em-eta9-phi11*/	4,86,1,7,86,2,5,163,3,6,164,3,9,
/* out0230_em-eta10-phi11*/	5,20,0,3,20,1,6,86,1,8,163,2,12,163,3,10,
/* out0231_em-eta11-phi11*/	8,20,1,8,20,2,2,20,4,2,21,0,6,21,1,16,110,0,2,114,0,10,163,2,4,
/* out0232_em-eta12-phi11*/	9,20,4,14,20,5,6,21,0,2,29,2,5,110,0,5,113,0,4,113,2,1,114,0,1,114,1,1,
/* out0233_em-eta13-phi11*/	7,28,5,2,29,0,1,29,2,3,29,4,6,29,5,13,109,0,1,113,0,9,
/* out0234_em-eta14-phi11*/	9,28,4,1,28,5,3,29,0,13,29,1,1,29,4,1,109,0,5,112,0,1,113,0,1,113,1,1,
/* out0235_em-eta15-phi11*/	6,4,0,1,28,4,2,29,0,1,29,1,13,109,0,2,112,0,6,
/* out0236_em-eta16-phi11*/	4,4,0,12,29,1,1,108,0,2,112,0,4,
/* out0237_em-eta17-phi11*/	4,4,0,2,4,1,9,108,0,4,111,2,1,
/* out0238_em-eta18-phi11*/	5,4,1,5,5,1,4,108,0,1,111,1,1,111,2,3,
/* out0239_em-eta19-phi11*/	1,5,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	1,172,0,16,
/* out0242_em-eta2-phi12*/	2,171,0,1,172,1,16,
/* out0243_em-eta3-phi12*/	8,128,1,7,128,2,1,129,1,1,129,2,2,130,0,15,130,2,9,171,0,15,171,1,3,
/* out0244_em-eta4-phi12*/	6,127,2,9,128,1,1,128,2,15,129,1,6,170,0,3,171,1,13,
/* out0245_em-eta5-phi12*/	6,126,0,2,127,0,5,127,1,16,127,2,4,170,0,13,170,1,5,
/* out0246_em-eta6-phi12*/	5,88,1,3,126,0,14,126,1,4,169,0,6,170,1,11,
/* out0247_em-eta7-phi12*/	5,87,1,4,87,2,9,126,1,5,169,0,10,169,1,7,
/* out0248_em-eta8-phi12*/	4,86,2,3,87,1,12,169,1,9,169,2,7,
/* out0249_em-eta9-phi12*/	4,86,0,6,86,2,6,168,0,6,169,2,9,
/* out0250_em-eta10-phi12*/	5,31,2,3,31,3,6,86,0,8,168,0,10,168,1,12,
/* out0251_em-eta11-phi12*/	7,31,2,13,31,3,4,31,4,8,31,5,9,110,0,2,110,1,8,168,1,4,
/* out0252_em-eta12-phi12*/	8,29,2,5,30,4,1,30,5,13,31,0,1,31,5,7,110,0,6,110,1,2,110,2,5,
/* out0253_em-eta13-phi12*/	9,28,2,1,28,3,1,29,2,3,29,3,12,29,4,7,109,0,1,109,1,5,110,0,1,110,2,4,
/* out0254_em-eta14-phi12*/	8,28,1,1,28,2,14,28,3,2,29,0,1,29,4,2,109,0,5,109,1,2,109,2,1,
/* out0255_em-eta15-phi12*/	8,28,0,1,28,1,14,28,2,1,29,1,1,37,5,1,108,1,1,109,0,2,109,2,5,
/* out0256_em-eta16-phi12*/	5,28,1,1,36,5,6,37,5,7,108,0,3,108,1,4,
/* out0257_em-eta17-phi12*/	4,36,4,3,36,5,8,108,0,4,108,2,1,
/* out0258_em-eta18-phi12*/	3,36,4,9,108,0,2,108,2,3,
/* out0259_em-eta19-phi12*/	1,36,4,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	1,172,3,16,
/* out0262_em-eta2-phi13*/	5,130,2,2,131,0,12,131,2,2,171,3,1,172,2,16,
/* out0263_em-eta3-phi13*/	10,90,1,1,129,0,3,129,2,13,130,0,1,130,2,5,131,0,2,131,1,5,131,2,14,171,2,3,171,3,15,
/* out0264_em-eta4-phi13*/	8,89,2,6,127,0,1,127,2,3,129,0,13,129,1,9,129,2,1,170,3,3,171,2,13,
/* out0265_em-eta5-phi13*/	6,88,2,6,89,1,3,89,2,7,127,0,10,170,2,5,170,3,13,
/* out0266_em-eta6-phi13*/	5,88,0,4,88,1,10,88,2,8,169,5,6,170,2,11,
/* out0267_em-eta7-phi13*/	7,87,0,5,87,2,7,88,0,2,88,1,3,99,1,1,169,4,7,169,5,10,
/* out0268_em-eta8-phi13*/	4,87,0,11,98,2,3,169,3,7,169,4,9,
/* out0269_em-eta9-phi13*/	5,86,0,1,98,1,1,98,2,11,168,3,6,169,3,9,
/* out0270_em-eta10-phi13*/	8,30,0,2,30,3,13,31,3,5,86,0,1,98,1,3,98,2,1,168,2,12,168,3,10,
/* out0271_em-eta11-phi13*/	10,30,0,1,30,1,1,30,2,16,30,3,3,31,0,6,31,3,1,31,4,8,107,0,10,110,1,4,168,2,4,
/* out0272_em-eta12-phi13*/	9,30,4,11,30,5,3,31,0,9,31,1,6,105,0,4,105,1,1,107,2,1,110,1,2,110,2,6,
/* out0273_em-eta13-phi13*/	8,28,3,8,29,3,4,30,4,3,38,5,6,39,5,3,105,0,5,109,1,5,110,2,1,
/* out0274_em-eta14-phi13*/	6,28,0,9,28,3,5,38,4,4,38,5,1,109,1,4,109,2,5,
/* out0275_em-eta15-phi13*/	6,28,0,6,37,2,9,37,5,1,103,0,2,108,1,1,109,2,5,
/* out0276_em-eta16-phi13*/	5,37,0,1,37,2,1,37,4,6,37,5,7,108,1,6,
/* out0277_em-eta17-phi13*/	5,36,5,2,37,0,9,37,4,1,108,1,1,108,2,4,
/* out0278_em-eta18-phi13*/	4,36,4,2,37,0,2,37,1,5,108,2,4,
/* out0279_em-eta19-phi13*/	2,36,4,1,37,1,3,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	1,177,0,16,
/* out0282_em-eta2-phi14*/	6,91,0,4,91,1,5,131,0,2,131,1,4,176,0,1,177,1,16,
/* out0283_em-eta3-phi14*/	8,90,0,4,90,1,4,90,2,16,91,0,1,91,1,10,131,1,7,176,0,15,176,1,3,
/* out0284_em-eta4-phi14*/	7,89,0,11,89,2,2,90,0,5,90,1,11,101,2,3,175,0,3,176,1,13,
/* out0285_em-eta5-phi14*/	7,88,2,1,89,0,5,89,1,13,89,2,1,100,2,6,175,0,13,175,1,5,
/* out0286_em-eta6-phi14*/	7,88,0,9,88,2,1,99,2,2,100,1,3,100,2,8,174,0,6,175,1,11,
/* out0287_em-eta7-phi14*/	6,88,0,1,99,0,1,99,1,6,99,2,11,174,0,10,174,1,7,
/* out0288_em-eta8-phi14*/	5,98,0,6,99,0,1,99,1,9,174,1,9,174,2,7,
/* out0289_em-eta9-phi14*/	5,98,0,7,98,1,4,98,2,1,173,0,6,174,2,9,
/* out0290_em-eta10-phi14*/	5,30,0,5,41,2,10,98,1,7,173,0,10,173,1,12,
/* out0291_em-eta11-phi14*/	7,30,0,8,30,1,13,41,2,5,41,5,8,107,0,6,107,2,13,173,1,4,
/* out0292_em-eta12-phi14*/	10,30,1,2,30,4,1,31,1,10,39,2,10,39,5,4,40,5,1,41,5,1,105,0,2,105,1,10,107,2,1,
/* out0293_em-eta13-phi14*/	6,38,5,5,39,0,5,39,4,6,39,5,9,105,0,5,105,2,6,
/* out0294_em-eta14-phi14*/	7,38,4,8,38,5,4,39,0,5,39,1,3,103,0,2,103,1,4,105,2,2,
/* out0295_em-eta15-phi14*/	5,37,2,6,37,3,5,38,4,4,39,1,2,103,0,7,
/* out0296_em-eta16-phi14*/	6,36,2,2,37,3,4,37,4,8,103,0,4,103,2,1,108,1,2,
/* out0297_em-eta17-phi14*/	6,36,2,8,37,0,2,37,4,1,102,1,2,108,1,1,108,2,3,
/* out0298_em-eta18-phi14*/	7,36,1,4,36,2,2,37,0,2,37,1,3,102,0,1,102,1,2,108,2,1,
/* out0299_em-eta19-phi14*/	2,36,1,2,37,1,5,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	1,177,3,16,
/* out0302_em-eta2-phi15*/	3,91,0,3,176,3,1,177,2,16,
/* out0303_em-eta3-phi15*/	8,90,0,4,91,0,8,91,1,1,102,0,7,102,1,6,102,2,16,176,2,3,176,3,15,
/* out0304_em-eta4-phi15*/	7,90,0,3,101,0,12,101,1,3,101,2,11,102,1,4,175,3,3,176,2,13,
/* out0305_em-eta5-phi15*/	7,100,0,11,100,2,1,101,1,11,101,2,2,110,1,1,175,2,5,175,3,13,
/* out0306_em-eta6-phi15*/	6,100,0,4,100,1,13,100,2,1,109,2,3,174,5,6,175,2,11,
/* out0307_em-eta7-phi15*/	6,99,0,9,99,2,3,109,1,5,109,2,1,174,4,7,174,5,10,
/* out0308_em-eta8-phi15*/	5,99,0,5,108,1,2,108,2,8,174,3,7,174,4,9,
/* out0309_em-eta9-phi15*/	7,40,3,1,41,3,1,98,0,3,98,1,1,108,1,9,173,3,6,174,3,9,
/* out0310_em-eta10-phi15*/	8,40,2,6,40,3,11,41,2,1,41,3,15,41,4,7,106,0,1,173,2,12,173,3,10,
/* out0311_em-eta11-phi15*/	10,40,2,1,40,5,7,41,0,9,41,4,9,41,5,7,106,0,7,106,1,1,106,2,11,107,2,1,173,2,4,
/* out0312_em-eta12-phi15*/	8,39,2,6,39,3,12,40,4,4,40,5,8,105,1,5,105,2,1,106,1,2,106,2,5,
/* out0313_em-eta13-phi15*/	7,38,2,9,38,3,2,39,0,1,39,3,2,39,4,10,104,1,4,105,2,7,
/* out0314_em-eta14-phi15*/	6,38,1,5,38,2,6,39,0,5,39,1,4,103,1,8,104,1,1,
/* out0315_em-eta15-phi15*/	8,13,2,1,36,3,1,37,3,5,38,1,3,39,1,7,103,0,1,103,1,2,103,2,4,
/* out0316_em-eta16-phi15*/	5,36,2,1,36,3,11,37,3,2,102,1,1,103,2,5,
/* out0317_em-eta17-phi15*/	5,36,0,4,36,1,1,36,2,3,36,3,3,102,1,5,
/* out0318_em-eta18-phi15*/	4,36,0,3,36,1,7,102,0,3,102,1,2,
/* out0319_em-eta19-phi15*/	6,8,3,3,8,5,1,9,3,2,9,5,2,36,1,2,102,0,2,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	1,182,0,16,
/* out0322_em-eta2-phi16*/	2,181,0,1,182,1,16,
/* out0323_em-eta3-phi16*/	8,102,0,9,102,1,5,111,0,4,111,2,2,112,0,4,112,1,14,181,0,15,181,1,3,
/* out0324_em-eta4-phi16*/	9,101,0,4,101,1,1,102,1,1,110,2,1,111,0,3,111,1,8,111,2,14,180,0,3,181,1,13,
/* out0325_em-eta5-phi16*/	6,101,1,1,110,0,4,110,1,7,110,2,14,180,0,13,180,1,5,
/* out0326_em-eta6-phi16*/	7,100,0,1,109,0,2,109,2,11,110,0,1,110,1,8,179,0,6,180,1,11,
/* out0327_em-eta7-phi16*/	5,109,0,7,109,1,10,109,2,1,179,0,10,179,1,7,
/* out0328_em-eta8-phi16*/	5,108,0,6,108,2,8,109,1,1,179,1,9,179,2,7,
/* out0329_em-eta9-phi16*/	4,108,0,7,108,1,5,178,0,6,179,2,9,
/* out0330_em-eta10-phi16*/	7,40,0,16,40,1,9,40,2,5,40,3,4,52,0,1,178,0,10,178,1,12,
/* out0331_em-eta11-phi16*/	8,40,1,5,40,2,4,40,4,3,41,0,7,41,1,14,106,0,8,106,1,8,178,1,4,
/* out0332_em-eta12-phi16*/	7,14,5,6,15,5,7,38,3,3,39,3,2,40,4,9,104,2,7,106,1,5,
/* out0333_em-eta13-phi16*/	8,14,4,2,14,5,3,38,0,7,38,2,1,38,3,11,104,0,1,104,1,7,104,2,3,
/* out0334_em-eta14-phi16*/	6,13,3,4,38,0,9,38,1,6,103,1,2,104,0,2,104,1,4,
/* out0335_em-eta15-phi16*/	5,13,2,11,13,3,4,38,1,2,98,1,3,103,2,4,
/* out0336_em-eta16-phi16*/	8,13,2,4,13,5,7,36,0,1,36,3,1,98,1,2,102,1,1,102,2,1,103,2,2,
/* out0337_em-eta17-phi16*/	6,8,0,1,12,5,1,13,5,4,36,0,6,102,1,2,102,2,3,
/* out0338_em-eta18-phi16*/	6,8,0,6,8,3,5,36,0,2,102,0,5,102,1,1,102,2,1,
/* out0339_em-eta19-phi16*/	6,8,2,1,8,3,6,8,5,5,9,3,9,9,5,9,102,0,3,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	1,182,3,16,
/* out0342_em-eta2-phi17*/	2,181,3,1,182,2,16,
/* out0343_em-eta3-phi17*/	5,111,0,3,112,0,12,112,1,2,181,2,3,181,3,15,
/* out0344_em-eta4-phi17*/	6,55,0,8,55,1,4,111,0,6,111,1,8,180,3,3,181,2,13,
/* out0345_em-eta5-phi17*/	8,54,0,1,54,1,2,55,0,8,55,2,4,110,0,9,110,2,1,180,2,5,180,3,13,
/* out0346_em-eta6-phi17*/	7,54,0,14,54,1,1,54,2,2,109,0,2,110,0,2,179,5,6,180,2,11,
/* out0347_em-eta7-phi17*/	6,53,1,10,54,0,1,54,2,2,109,0,5,179,4,7,179,5,10,
/* out0348_em-eta8-phi17*/	5,53,0,11,53,1,2,108,0,1,179,3,7,179,4,9,
/* out0349_em-eta9-phi17*/	6,52,0,6,52,1,4,53,0,1,108,0,2,178,3,6,179,3,9,
/* out0350_em-eta10-phi17*/	4,52,0,8,52,2,2,178,2,12,178,3,10,
/* out0351_em-eta11-phi17*/	10,15,2,16,15,3,4,15,5,1,40,1,2,41,1,2,52,0,1,52,2,2,101,0,9,101,2,7,178,2,4,
/* out0352_em-eta12-phi17*/	7,14,5,3,15,0,7,15,4,11,15,5,8,101,1,1,101,2,9,104,2,4,
/* out0353_em-eta13-phi17*/	6,14,4,11,14,5,4,15,0,5,15,1,3,104,0,8,104,2,2,
/* out0354_em-eta14-phi17*/	5,12,3,12,13,3,5,14,4,3,98,2,4,104,0,5,
/* out0355_em-eta15-phi17*/	5,12,2,4,13,3,3,13,4,10,98,1,4,98,2,3,
/* out0356_em-eta16-phi17*/	5,12,5,1,13,0,4,13,4,6,13,5,4,98,1,6,
/* out0357_em-eta17-phi17*/	5,8,0,2,12,5,10,13,5,1,98,1,1,102,2,5,
/* out0358_em-eta18-phi17*/	5,8,0,7,8,1,3,8,2,6,8,3,2,102,2,5,
/* out0359_em-eta19-phi17*/	7,8,2,5,8,5,8,9,0,4,9,3,5,9,5,5,102,0,2,102,2,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	1,187,0,16,
/* out0362_em-eta2-phi18*/	2,186,0,1,187,1,16,
/* out0363_em-eta3-phi18*/	6,64,0,1,64,1,2,65,0,11,65,2,3,186,0,15,186,1,3,
/* out0364_em-eta4-phi18*/	5,55,1,12,64,0,13,64,2,1,185,0,3,186,1,13,
/* out0365_em-eta5-phi18*/	6,54,1,4,55,2,12,63,0,9,63,1,1,185,0,13,185,1,5,
/* out0366_em-eta6-phi18*/	6,54,1,9,54,2,9,62,0,2,63,0,2,184,0,6,185,1,11,
/* out0367_em-eta7-phi18*/	6,53,1,4,53,2,6,54,2,3,62,0,5,184,0,10,184,1,7,
/* out0368_em-eta8-phi18*/	5,53,0,3,53,2,10,61,1,2,184,1,9,184,2,7,
/* out0369_em-eta9-phi18*/	5,52,1,10,53,0,1,61,0,2,183,0,6,184,2,9,
/* out0370_em-eta10-phi18*/	4,52,1,2,52,2,9,183,0,10,183,1,12,
/* out0371_em-eta11-phi18*/	9,14,3,8,15,3,12,15,4,1,26,5,2,27,5,2,52,2,2,101,0,7,101,1,7,183,1,4,
/* out0372_em-eta12-phi18*/	8,14,0,1,14,1,2,14,2,14,14,3,6,15,0,1,15,4,4,99,2,4,101,1,8,
/* out0373_em-eta13-phi18*/	6,14,1,9,14,2,2,15,0,3,15,1,10,99,1,8,99,2,2,
/* out0374_em-eta14-phi18*/	5,12,0,12,12,3,4,15,1,3,98,2,4,99,1,5,
/* out0375_em-eta15-phi18*/	5,12,1,3,12,2,12,13,0,2,98,0,4,98,2,4,
/* out0376_em-eta16-phi18*/	5,12,4,1,12,5,1,13,0,10,13,1,2,98,0,6,
/* out0377_em-eta17-phi18*/	5,8,1,2,12,4,8,12,5,3,98,0,1,128,1,4,
/* out0378_em-eta18-phi18*/	5,8,1,10,8,2,4,9,0,7,9,1,4,128,1,4,
/* out0379_em-eta19-phi18*/	6,8,4,5,8,5,2,9,0,5,9,1,1,128,0,2,128,1,1,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	1,187,3,16,
/* out0382_em-eta2-phi19*/	2,186,3,1,187,2,16,
/* out0383_em-eta3-phi19*/	7,64,1,6,65,0,5,65,2,13,75,0,5,75,1,9,186,2,3,186,3,15,
/* out0384_em-eta4-phi19*/	8,63,1,1,64,0,2,64,1,8,64,2,15,74,0,5,75,0,1,185,3,3,186,2,13,
/* out0385_em-eta5-phi19*/	6,63,0,4,63,1,14,63,2,7,74,0,1,185,2,5,185,3,13,
/* out0386_em-eta6-phi19*/	7,62,0,2,62,1,11,63,0,1,63,2,8,73,0,1,184,5,6,185,2,11,
/* out0387_em-eta7-phi19*/	5,62,0,7,62,1,2,62,2,10,184,4,7,184,5,10,
/* out0388_em-eta8-phi19*/	5,61,1,13,61,2,1,62,2,1,184,3,7,184,4,9,
/* out0389_em-eta9-phi19*/	3,61,0,11,183,3,6,184,3,9,
/* out0390_em-eta10-phi19*/	7,27,2,16,27,3,4,27,4,5,27,5,9,52,2,1,183,2,12,183,3,10,
/* out0391_em-eta11-phi19*/	10,14,3,1,26,4,3,26,5,14,27,0,7,27,4,4,27,5,5,100,0,10,100,1,1,100,2,8,183,2,4,
/* out0392_em-eta12-phi19*/	6,14,0,13,14,3,1,23,2,6,26,4,9,99,2,7,100,2,7,
/* out0393_em-eta13-phi19*/	7,14,0,2,14,1,5,23,2,4,23,5,14,99,0,7,99,1,1,99,2,3,
/* out0394_em-eta14-phi19*/	9,12,0,4,12,1,1,22,4,1,22,5,13,23,5,1,98,2,1,99,0,4,99,1,2,129,2,2,
/* out0395_em-eta15-phi19*/	5,12,1,12,13,1,3,22,4,2,98,0,3,129,1,4,
/* out0396_em-eta16-phi19*/	8,11,2,1,11,3,1,12,4,2,13,1,10,98,0,2,128,1,1,128,2,1,129,1,2,
/* out0397_em-eta17-phi19*/	5,8,1,1,11,2,6,12,4,5,128,1,4,128,2,1,
/* out0398_em-eta18-phi19*/	5,8,4,2,9,1,11,11,2,2,128,0,3,128,1,2,
/* out0399_em-eta19-phi19*/	2,8,4,6,128,0,3,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	1,192,0,16,
/* out0402_em-eta2-phi20*/	3,85,0,3,191,0,1,192,1,16,
/* out0403_em-eta3-phi20*/	8,75,0,6,75,1,7,75,2,16,84,1,4,85,0,8,85,2,1,191,0,15,191,1,3,
/* out0404_em-eta4-phi20*/	8,74,0,6,74,1,15,74,2,5,75,0,4,84,0,2,84,1,1,190,0,3,191,1,13,
/* out0405_em-eta5-phi20*/	7,63,2,1,73,0,3,73,1,9,74,0,4,74,2,9,190,0,13,190,1,5,
/* out0406_em-eta6-phi20*/	6,62,1,2,73,0,12,73,1,1,73,2,6,189,0,6,190,1,11,
/* out0407_em-eta7-phi20*/	6,62,1,1,62,2,5,72,0,9,72,1,3,189,0,10,189,1,7,
/* out0408_em-eta8-phi20*/	5,61,1,1,61,2,9,72,0,5,189,1,9,189,2,7,
/* out0409_em-eta9-phi20*/	7,26,3,1,27,3,1,61,0,3,61,2,6,71,0,3,188,0,6,189,2,9,
/* out0410_em-eta10-phi20*/	9,26,0,1,26,2,7,26,3,15,27,3,11,27,4,6,71,0,1,100,0,1,188,0,10,188,1,12,
/* out0411_em-eta11-phi20*/	9,26,1,7,26,2,9,27,0,9,27,1,7,27,4,1,100,0,5,100,1,10,131,1,1,188,1,4,
/* out0412_em-eta12-phi20*/	8,23,2,5,23,3,12,26,4,4,27,1,8,100,1,5,100,2,1,130,1,1,130,2,5,
/* out0413_em-eta13-phi20*/	8,22,2,3,23,0,2,23,2,1,23,3,2,23,4,16,23,5,1,99,0,4,130,1,7,
/* out0414_em-eta14-phi20*/	6,22,4,3,22,5,3,23,0,11,23,1,3,99,0,1,129,2,8,
/* out0415_em-eta15-phi20*/	8,10,3,5,11,3,1,13,1,1,22,4,10,23,1,1,129,0,1,129,1,4,129,2,2,
/* out0416_em-eta16-phi20*/	5,10,3,2,11,3,11,11,4,1,128,2,1,129,1,5,
/* out0417_em-eta17-phi20*/	5,11,2,4,11,3,3,11,4,3,11,5,1,128,2,6,
/* out0418_em-eta18-phi20*/	4,11,2,3,11,5,7,128,0,5,128,2,2,
/* out0419_em-eta19-phi20*/	3,8,4,3,11,5,2,128,0,2,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	1,192,3,16,
/* out0422_em-eta2-phi21*/	6,85,0,4,85,2,5,125,0,3,125,2,4,191,3,1,192,2,16,
/* out0423_em-eta3-phi21*/	8,84,0,1,84,1,11,84,2,12,85,0,1,85,2,10,125,2,9,191,2,3,191,3,15,
/* out0424_em-eta4-phi21*/	8,74,1,1,74,2,2,83,0,3,83,1,10,84,0,13,84,2,3,190,3,3,191,2,13,
/* out0425_em-eta5-phi21*/	7,73,1,6,82,1,1,83,0,13,83,1,1,83,2,5,190,2,5,190,3,13,
/* out0426_em-eta6-phi21*/	6,72,1,2,73,2,10,82,0,9,82,1,1,189,5,6,190,2,11,
/* out0427_em-eta7-phi21*/	6,72,0,1,72,1,11,72,2,6,82,0,1,189,4,7,189,5,10,
/* out0428_em-eta8-phi21*/	5,71,1,6,72,0,1,72,2,9,189,3,7,189,4,9,
/* out0429_em-eta9-phi21*/	5,71,0,8,71,1,3,71,2,1,188,3,6,189,3,9,
/* out0430_em-eta10-phi21*/	6,25,2,5,26,0,10,71,0,4,71,2,3,188,2,12,188,3,10,
/* out0431_em-eta11-phi21*/	7,25,2,8,25,5,13,26,0,5,26,1,8,131,0,6,131,1,13,188,2,4,
/* out0432_em-eta12-phi21*/	11,22,0,1,22,3,11,23,3,2,24,4,1,24,5,10,25,5,2,26,1,1,27,1,1,130,0,2,130,2,10,131,1,1,
/* out0433_em-eta13-phi21*/	6,22,0,6,22,1,3,22,2,10,22,3,5,130,0,5,130,1,6,
/* out0434_em-eta14-phi21*/	7,22,1,8,22,2,3,23,0,3,23,1,7,129,0,2,129,2,4,130,1,2,
/* out0435_em-eta15-phi21*/	4,10,0,6,10,3,5,23,1,5,129,0,7,
/* out0436_em-eta16-phi21*/	6,10,2,8,10,3,4,11,4,2,95,2,2,129,0,4,129,1,1,
/* out0437_em-eta17-phi21*/	6,10,2,1,11,0,2,11,4,8,95,1,3,95,2,1,128,2,2,
/* out0438_em-eta18-phi21*/	7,10,5,3,11,0,2,11,4,2,11,5,4,95,1,1,128,0,1,128,2,3,
/* out0439_em-eta19-phi21*/	2,10,5,5,11,5,2,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	1,197,0,16,
/* out0442_em-eta2-phi22*/	5,124,0,2,125,0,12,125,1,2,196,0,1,197,1,16,
/* out0443_em-eta3-phi22*/	10,84,2,1,123,0,3,123,1,13,124,0,5,124,2,1,125,0,1,125,1,14,125,2,3,196,0,15,196,1,3,
/* out0444_em-eta4-phi22*/	9,83,1,5,83,2,1,122,0,1,122,1,3,123,0,13,123,1,1,123,2,9,195,0,3,196,1,13,
/* out0445_em-eta5-phi22*/	5,82,1,6,83,2,10,122,0,10,195,0,13,195,1,5,
/* out0446_em-eta6-phi22*/	5,82,0,4,82,1,8,82,2,10,194,0,6,195,1,11,
/* out0447_em-eta7-phi22*/	7,72,2,1,81,0,5,81,1,7,82,0,2,82,2,3,194,0,10,194,1,7,
/* out0448_em-eta8-phi22*/	4,71,1,3,81,0,11,194,1,9,194,2,7,
/* out0449_em-eta9-phi22*/	4,71,1,4,71,2,8,193,0,6,194,2,9,
/* out0450_em-eta10-phi22*/	6,24,3,5,25,2,2,25,3,13,71,2,4,193,0,10,193,1,12,
/* out0451_em-eta11-phi22*/	10,24,2,8,24,3,1,25,0,6,25,2,1,25,3,3,25,4,16,25,5,1,97,2,4,131,0,10,193,1,4,
/* out0452_em-eta12-phi22*/	9,24,4,11,24,5,6,25,0,9,25,1,3,97,1,6,97,2,2,130,0,4,130,2,1,131,1,1,
/* out0453_em-eta13-phi22*/	5,22,0,9,24,4,3,96,2,5,97,1,1,130,0,5,
/* out0454_em-eta14-phi22*/	3,22,1,5,96,1,5,96,2,4,
/* out0455_em-eta15-phi22*/	5,10,0,9,10,1,1,95,2,1,96,1,5,129,0,2,
/* out0456_em-eta16-phi22*/	5,10,0,1,10,1,7,10,2,6,11,0,1,95,2,6,
/* out0457_em-eta17-phi22*/	5,10,2,1,11,0,9,11,1,2,95,1,4,95,2,1,
/* out0458_em-eta18-phi22*/	4,10,4,2,10,5,5,11,0,2,95,1,4,
/* out0459_em-eta19-phi22*/	2,10,4,1,10,5,3,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	1,197,3,16,
/* out0462_em-eta2-phi23*/	2,196,3,1,197,2,16,
/* out0463_em-eta3-phi23*/	6,123,1,2,123,2,1,124,0,9,124,2,15,196,2,3,196,3,15,
/* out0464_em-eta4-phi23*/	4,122,1,9,123,2,6,195,3,3,196,2,13,
/* out0465_em-eta5-phi23*/	5,122,0,5,122,1,4,122,2,16,195,2,5,195,3,13,
/* out0466_em-eta6-phi23*/	3,82,2,3,194,5,6,195,2,11,
/* out0467_em-eta7-phi23*/	4,81,1,9,81,2,4,194,4,7,194,5,10,
/* out0468_em-eta8-phi23*/	3,81,2,12,194,3,7,194,4,9,
/* out0469_em-eta9-phi23*/	2,193,3,6,194,3,9,
/* out0470_em-eta10-phi23*/	4,24,0,3,24,3,6,193,2,12,193,3,10,
/* out0471_em-eta11-phi23*/	7,24,0,13,24,1,9,24,2,8,24,3,4,97,0,9,97,2,8,193,2,4,
/* out0472_em-eta12-phi23*/	7,24,1,7,24,4,1,25,0,1,25,1,13,97,0,6,97,1,5,97,2,2,
/* out0473_em-eta13-phi23*/	4,96,0,2,96,2,5,97,0,1,97,1,4,
/* out0474_em-eta14-phi23*/	3,96,0,12,96,1,1,96,2,2,
/* out0475_em-eta15-phi23*/	5,10,1,1,95,0,1,95,2,1,96,0,2,96,1,5,
/* out0476_em-eta16-phi23*/	4,10,1,7,11,1,6,95,0,3,95,2,4,
/* out0477_em-eta17-phi23*/	4,10,4,3,11,1,8,95,0,5,95,1,1,
/* out0478_em-eta18-phi23*/	3,10,4,9,95,0,2,95,1,3,
/* out0479_em-eta19-phi23*/	2,10,4,1,95,0,5
};