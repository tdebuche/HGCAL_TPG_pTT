parameter integer matrixH [0:6372] = {
/* num inputs = 170(in0-in169) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 10 */
//* total number of input in adders 1964 */

/* out0000_had-eta0-phi0*/	1, 125, 0, 6, 
/* out0001_had-eta1-phi0*/	2, 124, 0, 3, 125, 0, 10, 
/* out0002_had-eta2-phi0*/	2, 124, 0, 13, 124, 1, 5, 
/* out0003_had-eta3-phi0*/	4, 36, 1, 6, 36, 2, 11, 123, 0, 6, 124, 1, 11, 
/* out0004_had-eta4-phi0*/	6, 27, 2, 12, 35, 1, 2, 35, 2, 9, 36, 1, 4, 123, 0, 10, 123, 1, 7, 
/* out0005_had-eta5-phi0*/	7, 27, 0, 15, 27, 1, 2, 27, 2, 4, 34, 2, 4, 35, 1, 6, 122, 0, 8, 123, 1, 9, 
/* out0006_had-eta6-phi0*/	8, 26, 0, 8, 26, 2, 5, 27, 0, 1, 27, 1, 14, 34, 1, 5, 34, 2, 3, 122, 0, 8, 122, 1, 16, 
/* out0007_had-eta7-phi0*/	6, 25, 2, 13, 26, 0, 8, 26, 1, 16, 26, 2, 11, 33, 1, 2, 33, 2, 4, 
/* out0008_had-eta8-phi0*/	4, 25, 0, 12, 25, 1, 12, 25, 2, 3, 33, 1, 2, 
/* out0009_had-eta9-phi0*/	6, 24, 0, 1, 24, 2, 14, 25, 0, 4, 25, 1, 4, 32, 1, 1, 32, 2, 2, 
/* out0010_had-eta10-phi0*/	3, 24, 0, 9, 24, 1, 12, 24, 2, 2, 
/* out0011_had-eta11-phi0*/	6, 3, 8, 16, 3, 9, 3, 9, 5, 1, 9, 11, 2, 24, 0, 4, 24, 1, 4, 
/* out0012_had-eta12-phi0*/	5, 3, 2, 4, 3, 3, 13, 3, 9, 13, 3, 10, 4, 9, 5, 1, 
/* out0013_had-eta13-phi0*/	7, 3, 0, 1, 3, 1, 7, 3, 2, 12, 3, 3, 1, 3, 6, 16, 3, 7, 1, 3, 10, 12, 
/* out0014_had-eta14-phi0*/	6, 1, 3, 1, 1, 8, 16, 1, 9, 9, 3, 1, 4, 3, 4, 16, 3, 7, 15, 
/* out0015_had-eta15-phi0*/	4, 1, 2, 3, 1, 3, 6, 1, 9, 7, 1, 10, 4, 
/* out0016_had-eta16-phi0*/	3, 1, 2, 12, 1, 6, 13, 1, 10, 12, 
/* out0017_had-eta17-phi0*/	4, 1, 1, 3, 1, 2, 1, 1, 6, 3, 1, 7, 7, 
/* out0018_had-eta18-phi0*/	4, 0, 3, 16, 0, 4, 6, 1, 4, 16, 1, 7, 6, 
/* out0019_had-eta19-phi0*/	4, 0, 1, 5, 0, 2, 1, 0, 4, 6, 0, 5, 16, 
/* out0020_had-eta0-phi1*/	1, 125, 1, 6, 
/* out0021_had-eta1-phi1*/	2, 124, 3, 3, 125, 1, 10, 
/* out0022_had-eta2-phi1*/	2, 124, 2, 5, 124, 3, 13, 
/* out0023_had-eta3-phi1*/	7, 36, 0, 15, 36, 1, 2, 36, 2, 5, 46, 2, 6, 47, 1, 12, 123, 3, 6, 124, 2, 11, 
/* out0024_had-eta4-phi1*/	10, 35, 0, 12, 35, 1, 1, 35, 2, 7, 36, 0, 1, 36, 1, 4, 45, 2, 1, 46, 1, 7, 46, 2, 3, 123, 2, 7, 123, 3, 10, 
/* out0025_had-eta5-phi1*/	8, 34, 0, 5, 34, 2, 7, 35, 0, 4, 35, 1, 7, 45, 1, 3, 45, 2, 3, 122, 3, 8, 123, 2, 9, 
/* out0026_had-eta6-phi1*/	6, 33, 2, 2, 34, 0, 9, 34, 1, 11, 34, 2, 2, 122, 2, 16, 122, 3, 8, 
/* out0027_had-eta7-phi1*/	3, 33, 0, 7, 33, 1, 3, 33, 2, 10, 
/* out0028_had-eta8-phi1*/	3, 32, 2, 6, 33, 0, 1, 33, 1, 9, 
/* out0029_had-eta9-phi1*/	3, 32, 0, 1, 32, 1, 5, 32, 2, 7, 
/* out0030_had-eta10-phi1*/	4, 9, 8, 11, 9, 9, 2, 24, 0, 2, 32, 1, 7, 
/* out0031_had-eta11-phi1*/	6, 9, 5, 3, 9, 6, 4, 9, 8, 5, 9, 9, 1, 9, 10, 9, 9, 11, 14, 
/* out0032_had-eta12-phi1*/	5, 3, 0, 5, 3, 3, 2, 9, 4, 11, 9, 5, 11, 9, 6, 3, 
/* out0033_had-eta13-phi1*/	5, 3, 0, 10, 3, 1, 3, 8, 8, 10, 8, 11, 3, 9, 4, 1, 
/* out0034_had-eta14-phi1*/	4, 1, 3, 1, 3, 1, 2, 8, 5, 8, 8, 11, 12, 
/* out0035_had-eta15-phi1*/	4, 1, 0, 3, 1, 3, 7, 8, 4, 3, 8, 5, 5, 
/* out0036_had-eta16-phi1*/	3, 1, 0, 11, 1, 1, 3, 1, 3, 1, 
/* out0037_had-eta17-phi1*/	5, 1, 0, 1, 1, 1, 9, 1, 7, 2, 2, 8, 1, 2, 11, 3, 
/* out0038_had-eta18-phi1*/	6, 0, 2, 4, 0, 4, 2, 1, 1, 1, 1, 7, 1, 2, 5, 3, 2, 11, 2, 
/* out0039_had-eta19-phi1*/	4, 0, 0, 5, 0, 1, 11, 0, 2, 10, 0, 4, 2, 
/* out0040_had-eta0-phi2*/	1, 129, 0, 6, 
/* out0041_had-eta1-phi2*/	2, 128, 0, 3, 129, 0, 10, 
/* out0042_had-eta2-phi2*/	4, 47, 0, 2, 58, 2, 2, 128, 0, 13, 128, 1, 5, 
/* out0043_had-eta3-phi2*/	8, 46, 0, 7, 46, 2, 6, 47, 0, 14, 47, 1, 4, 58, 1, 9, 58, 2, 10, 127, 0, 6, 128, 1, 11, 
/* out0044_had-eta4-phi2*/	9, 45, 0, 3, 45, 2, 6, 46, 0, 9, 46, 1, 9, 46, 2, 1, 57, 1, 2, 57, 2, 5, 127, 0, 10, 127, 1, 7, 
/* out0045_had-eta5-phi2*/	6, 44, 2, 1, 45, 0, 10, 45, 1, 13, 45, 2, 6, 126, 0, 8, 127, 1, 9, 
/* out0046_had-eta6-phi2*/	6, 34, 0, 2, 44, 0, 3, 44, 1, 5, 44, 2, 15, 126, 0, 8, 126, 1, 16, 
/* out0047_had-eta7-phi2*/	3, 33, 0, 6, 43, 2, 6, 44, 1, 8, 
/* out0048_had-eta8-phi2*/	5, 32, 0, 3, 32, 2, 1, 33, 0, 2, 43, 1, 6, 43, 2, 5, 
/* out0049_had-eta9-phi2*/	3, 32, 0, 11, 42, 2, 2, 43, 1, 1, 
/* out0050_had-eta10-phi2*/	6, 9, 3, 9, 9, 9, 11, 32, 0, 1, 32, 1, 3, 42, 1, 1, 42, 2, 1, 
/* out0051_had-eta11-phi2*/	7, 9, 0, 2, 9, 1, 3, 9, 2, 15, 9, 3, 7, 9, 6, 3, 9, 9, 2, 9, 10, 7, 
/* out0052_had-eta12-phi2*/	6, 8, 9, 2, 9, 1, 4, 9, 2, 1, 9, 4, 4, 9, 6, 6, 9, 7, 15, 
/* out0053_had-eta13-phi2*/	5, 8, 2, 1, 8, 8, 6, 8, 9, 12, 8, 10, 7, 8, 11, 1, 
/* out0054_had-eta14-phi2*/	4, 8, 2, 2, 8, 5, 1, 8, 6, 11, 8, 10, 9, 
/* out0055_had-eta15-phi2*/	4, 8, 4, 11, 8, 5, 2, 8, 6, 2, 8, 7, 3, 
/* out0056_had-eta16-phi2*/	3, 1, 0, 1, 2, 8, 12, 8, 4, 2, 
/* out0057_had-eta17-phi2*/	3, 2, 8, 2, 2, 10, 2, 2, 11, 9, 
/* out0058_had-eta18-phi2*/	4, 2, 5, 7, 2, 6, 1, 2, 10, 1, 2, 11, 2, 
/* out0059_had-eta19-phi2*/	4, 0, 0, 11, 0, 2, 1, 2, 4, 4, 2, 5, 4, 
/* out0060_had-eta0-phi3*/	1, 129, 1, 6, 
/* out0061_had-eta1-phi3*/	2, 128, 3, 3, 129, 1, 10, 
/* out0062_had-eta2-phi3*/	4, 58, 0, 2, 58, 2, 2, 128, 2, 5, 128, 3, 13, 
/* out0063_had-eta3-phi3*/	9, 57, 0, 1, 57, 2, 3, 58, 0, 14, 58, 1, 7, 58, 2, 2, 100, 1, 4, 100, 2, 10, 127, 3, 6, 128, 2, 11, 
/* out0064_had-eta4-phi3*/	6, 57, 0, 14, 57, 1, 13, 57, 2, 8, 100, 1, 1, 127, 2, 7, 127, 3, 10, 
/* out0065_had-eta5-phi3*/	7, 45, 0, 3, 56, 0, 3, 56, 1, 6, 56, 2, 16, 57, 1, 1, 126, 3, 8, 127, 2, 9, 
/* out0066_had-eta6-phi3*/	5, 44, 0, 12, 55, 2, 6, 56, 1, 6, 126, 2, 16, 126, 3, 8, 
/* out0067_had-eta7-phi3*/	6, 43, 0, 6, 43, 2, 4, 44, 0, 1, 44, 1, 3, 55, 1, 4, 55, 2, 2, 
/* out0068_had-eta8-phi3*/	3, 43, 0, 8, 43, 1, 7, 43, 2, 1, 
/* out0069_had-eta9-phi3*/	3, 42, 0, 1, 42, 2, 11, 43, 1, 2, 
/* out0070_had-eta10-phi3*/	2, 42, 1, 9, 42, 2, 2, 
/* out0071_had-eta11-phi3*/	5, 9, 0, 14, 9, 1, 2, 10, 8, 13, 10, 11, 2, 42, 1, 2, 
/* out0072_had-eta12-phi3*/	6, 8, 3, 1, 8, 9, 1, 9, 1, 7, 9, 7, 1, 10, 5, 8, 10, 11, 14, 
/* out0073_had-eta13-phi3*/	6, 8, 0, 4, 8, 2, 3, 8, 3, 15, 8, 9, 1, 10, 4, 1, 10, 5, 3, 
/* out0074_had-eta14-phi3*/	4, 8, 0, 3, 8, 1, 7, 8, 2, 10, 8, 6, 2, 
/* out0075_had-eta15-phi3*/	4, 2, 9, 2, 8, 1, 3, 8, 6, 1, 8, 7, 13, 
/* out0076_had-eta16-phi3*/	3, 2, 8, 1, 2, 9, 12, 2, 10, 2, 
/* out0077_had-eta17-phi3*/	3, 2, 2, 2, 2, 6, 1, 2, 10, 11, 
/* out0078_had-eta18-phi3*/	2, 2, 5, 1, 2, 6, 10, 
/* out0079_had-eta19-phi3*/	3, 2, 4, 7, 2, 5, 1, 2, 7, 1, 
/* out0080_had-eta0-phi4*/	1, 133, 0, 6, 
/* out0081_had-eta1-phi4*/	2, 132, 0, 3, 133, 0, 10, 
/* out0082_had-eta2-phi4*/	5, 102, 0, 1, 102, 1, 5, 102, 2, 16, 132, 0, 13, 132, 1, 5, 
/* out0083_had-eta3-phi4*/	8, 100, 0, 16, 100, 1, 8, 100, 2, 6, 101, 1, 1, 101, 2, 5, 102, 1, 6, 131, 0, 6, 132, 1, 11, 
/* out0084_had-eta4-phi4*/	7, 57, 0, 1, 99, 0, 8, 99, 1, 8, 99, 2, 16, 100, 1, 3, 131, 0, 10, 131, 1, 7, 
/* out0085_had-eta5-phi4*/	6, 56, 0, 13, 56, 1, 1, 98, 2, 9, 99, 1, 7, 130, 0, 8, 131, 1, 9, 
/* out0086_had-eta6-phi4*/	7, 55, 0, 9, 55, 2, 7, 56, 1, 3, 98, 1, 4, 98, 2, 1, 130, 0, 8, 130, 1, 16, 
/* out0087_had-eta7-phi4*/	4, 54, 2, 3, 55, 0, 3, 55, 1, 12, 55, 2, 1, 
/* out0088_had-eta8-phi4*/	3, 43, 0, 2, 54, 1, 3, 54, 2, 11, 
/* out0089_had-eta9-phi4*/	2, 42, 0, 9, 54, 1, 5, 
/* out0090_had-eta10-phi4*/	4, 10, 9, 1, 42, 0, 6, 42, 1, 4, 64, 2, 1, 
/* out0091_had-eta11-phi4*/	5, 10, 2, 4, 10, 3, 6, 10, 8, 3, 10, 9, 15, 10, 10, 8, 
/* out0092_had-eta12-phi4*/	5, 10, 2, 4, 10, 5, 3, 10, 6, 15, 10, 7, 1, 10, 10, 8, 
/* out0093_had-eta13-phi4*/	5, 8, 0, 4, 10, 4, 14, 10, 5, 2, 10, 7, 2, 14, 8, 3, 
/* out0094_had-eta14-phi4*/	4, 8, 0, 5, 8, 1, 3, 14, 8, 7, 14, 11, 5, 
/* out0095_had-eta15-phi4*/	5, 2, 3, 1, 2, 9, 1, 8, 1, 3, 14, 5, 5, 14, 11, 7, 
/* out0096_had-eta16-phi4*/	3, 2, 2, 1, 2, 3, 13, 2, 9, 1, 
/* out0097_had-eta17-phi4*/	3, 2, 1, 1, 2, 2, 10, 2, 3, 2, 
/* out0098_had-eta18-phi4*/	4, 2, 1, 1, 2, 2, 3, 2, 6, 4, 2, 7, 2, 
/* out0099_had-eta19-phi4*/	2, 2, 4, 5, 2, 7, 8, 
/* out0100_had-eta0-phi5*/	1, 133, 1, 6, 
/* out0101_had-eta1-phi5*/	2, 132, 3, 3, 133, 1, 10, 
/* out0102_had-eta2-phi5*/	4, 102, 0, 14, 102, 1, 2, 132, 2, 5, 132, 3, 13, 
/* out0103_had-eta3-phi5*/	7, 101, 0, 16, 101, 1, 7, 101, 2, 11, 102, 0, 1, 102, 1, 3, 131, 3, 6, 132, 2, 11, 
/* out0104_had-eta4-phi5*/	6, 99, 0, 8, 101, 1, 8, 110, 1, 2, 110, 2, 16, 131, 2, 7, 131, 3, 10, 
/* out0105_had-eta5-phi5*/	7, 98, 0, 15, 98, 1, 1, 98, 2, 6, 99, 1, 1, 110, 1, 5, 130, 3, 8, 131, 2, 9, 
/* out0106_had-eta6-phi5*/	6, 55, 0, 2, 98, 0, 1, 98, 1, 11, 108, 2, 10, 130, 2, 16, 130, 3, 8, 
/* out0107_had-eta7-phi5*/	5, 54, 0, 3, 54, 2, 1, 55, 0, 2, 108, 1, 8, 108, 2, 6, 
/* out0108_had-eta8-phi5*/	3, 54, 0, 13, 54, 1, 3, 54, 2, 1, 
/* out0109_had-eta9-phi5*/	2, 54, 1, 5, 64, 2, 8, 
/* out0110_had-eta10-phi5*/	2, 64, 1, 5, 64, 2, 7, 
/* out0111_had-eta11-phi5*/	4, 10, 0, 13, 10, 2, 2, 10, 3, 10, 64, 1, 3, 
/* out0112_had-eta12-phi5*/	5, 10, 0, 3, 10, 1, 16, 10, 2, 6, 10, 6, 1, 10, 7, 5, 
/* out0113_had-eta13-phi5*/	4, 10, 4, 1, 10, 7, 8, 14, 8, 3, 14, 9, 12, 
/* out0114_had-eta14-phi5*/	4, 14, 8, 3, 14, 9, 3, 14, 10, 14, 14, 11, 3, 
/* out0115_had-eta15-phi5*/	4, 14, 5, 9, 14, 6, 7, 14, 10, 1, 14, 11, 1, 
/* out0116_had-eta16-phi5*/	3, 2, 0, 6, 14, 4, 7, 14, 5, 2, 
/* out0117_had-eta17-phi5*/	2, 2, 0, 10, 2, 1, 3, 
/* out0118_had-eta18-phi5*/	1, 2, 1, 10, 
/* out0119_had-eta19-phi5*/	2, 2, 1, 1, 2, 7, 5, 
/* out0120_had-eta0-phi6*/	1, 137, 0, 6, 
/* out0121_had-eta1-phi6*/	2, 136, 0, 3, 137, 0, 10, 
/* out0122_had-eta2-phi6*/	4, 114, 1, 1, 114, 2, 14, 136, 0, 13, 136, 1, 5, 
/* out0123_had-eta3-phi6*/	7, 112, 0, 11, 112, 1, 7, 112, 2, 16, 114, 1, 3, 114, 2, 1, 135, 0, 6, 136, 1, 11, 
/* out0124_had-eta4-phi6*/	6, 110, 0, 16, 110, 1, 3, 111, 2, 8, 112, 1, 8, 135, 0, 10, 135, 1, 7, 
/* out0125_had-eta5-phi6*/	7, 109, 0, 6, 109, 1, 1, 109, 2, 15, 110, 1, 6, 111, 1, 1, 134, 0, 8, 135, 1, 9, 
/* out0126_had-eta6-phi6*/	6, 66, 2, 2, 108, 0, 10, 109, 1, 11, 109, 2, 1, 134, 0, 8, 134, 1, 16, 
/* out0127_had-eta7-phi6*/	5, 65, 0, 1, 65, 2, 3, 66, 2, 2, 108, 0, 6, 108, 1, 8, 
/* out0128_had-eta8-phi6*/	3, 65, 0, 1, 65, 1, 3, 65, 2, 13, 
/* out0129_had-eta9-phi6*/	2, 64, 0, 8, 65, 1, 5, 
/* out0130_had-eta10-phi6*/	2, 64, 0, 7, 64, 1, 5, 
/* out0131_had-eta11-phi6*/	4, 15, 8, 13, 15, 9, 10, 15, 10, 2, 64, 1, 3, 
/* out0132_had-eta12-phi6*/	5, 15, 5, 5, 15, 6, 1, 15, 8, 3, 15, 10, 6, 15, 11, 16, 
/* out0133_had-eta13-phi6*/	5, 14, 0, 2, 14, 3, 13, 14, 9, 1, 15, 4, 1, 15, 5, 8, 
/* out0134_had-eta14-phi6*/	6, 14, 0, 2, 14, 1, 2, 14, 2, 15, 14, 3, 3, 14, 6, 1, 14, 10, 1, 
/* out0135_had-eta15-phi6*/	5, 14, 1, 1, 14, 2, 1, 14, 4, 1, 14, 6, 8, 14, 7, 8, 
/* out0136_had-eta16-phi6*/	3, 14, 4, 8, 14, 7, 1, 18, 8, 6, 
/* out0137_had-eta17-phi6*/	2, 18, 8, 10, 18, 11, 3, 
/* out0138_had-eta18-phi6*/	1, 18, 11, 10, 
/* out0139_had-eta19-phi6*/	2, 18, 5, 5, 18, 11, 1, 
/* out0140_had-eta0-phi7*/	1, 137, 1, 6, 
/* out0141_had-eta1-phi7*/	2, 136, 3, 3, 137, 1, 10, 
/* out0142_had-eta2-phi7*/	5, 114, 0, 16, 114, 1, 6, 114, 2, 1, 136, 2, 5, 136, 3, 13, 
/* out0143_had-eta3-phi7*/	8, 112, 0, 5, 112, 1, 1, 113, 0, 6, 113, 1, 8, 113, 2, 16, 114, 1, 6, 135, 3, 6, 136, 2, 11, 
/* out0144_had-eta4-phi7*/	7, 68, 2, 1, 111, 0, 16, 111, 1, 8, 111, 2, 8, 113, 1, 3, 135, 2, 7, 135, 3, 10, 
/* out0145_had-eta5-phi7*/	6, 67, 1, 1, 67, 2, 13, 109, 0, 9, 111, 1, 7, 134, 3, 8, 135, 2, 9, 
/* out0146_had-eta6-phi7*/	7, 66, 0, 7, 66, 2, 9, 67, 1, 3, 109, 0, 1, 109, 1, 4, 134, 2, 16, 134, 3, 8, 
/* out0147_had-eta7-phi7*/	4, 65, 0, 3, 66, 0, 1, 66, 1, 12, 66, 2, 3, 
/* out0148_had-eta8-phi7*/	3, 65, 0, 11, 65, 1, 3, 77, 2, 2, 
/* out0149_had-eta9-phi7*/	2, 65, 1, 5, 76, 2, 9, 
/* out0150_had-eta10-phi7*/	4, 15, 3, 1, 64, 0, 1, 76, 1, 4, 76, 2, 6, 
/* out0151_had-eta11-phi7*/	5, 15, 0, 3, 15, 2, 8, 15, 3, 15, 15, 9, 6, 15, 10, 4, 
/* out0152_had-eta12-phi7*/	5, 15, 2, 8, 15, 5, 1, 15, 6, 15, 15, 7, 3, 15, 10, 4, 
/* out0153_had-eta13-phi7*/	5, 14, 0, 4, 15, 4, 14, 15, 5, 2, 15, 7, 2, 19, 8, 4, 
/* out0154_had-eta14-phi7*/	4, 14, 0, 8, 14, 1, 6, 19, 8, 5, 19, 11, 3, 
/* out0155_had-eta15-phi7*/	5, 14, 1, 7, 14, 7, 6, 18, 3, 1, 18, 9, 1, 19, 11, 3, 
/* out0156_had-eta16-phi7*/	4, 14, 7, 1, 18, 3, 1, 18, 9, 13, 18, 10, 1, 
/* out0157_had-eta17-phi7*/	3, 18, 9, 2, 18, 10, 10, 18, 11, 1, 
/* out0158_had-eta18-phi7*/	4, 18, 5, 2, 18, 6, 4, 18, 10, 3, 18, 11, 1, 
/* out0159_had-eta19-phi7*/	2, 18, 4, 5, 18, 5, 8, 
/* out0160_had-eta0-phi8*/	1, 141, 0, 6, 
/* out0161_had-eta1-phi8*/	2, 140, 0, 3, 141, 0, 10, 
/* out0162_had-eta2-phi8*/	4, 69, 0, 2, 69, 2, 2, 140, 0, 13, 140, 1, 5, 
/* out0163_had-eta3-phi8*/	9, 68, 0, 3, 68, 2, 1, 69, 0, 2, 69, 1, 7, 69, 2, 14, 113, 0, 10, 113, 1, 4, 139, 0, 6, 140, 1, 11, 
/* out0164_had-eta4-phi8*/	6, 68, 0, 8, 68, 1, 13, 68, 2, 14, 113, 1, 1, 139, 0, 10, 139, 1, 7, 
/* out0165_had-eta5-phi8*/	7, 67, 0, 16, 67, 1, 6, 67, 2, 3, 68, 1, 1, 79, 2, 3, 138, 0, 8, 139, 1, 9, 
/* out0166_had-eta6-phi8*/	5, 66, 0, 6, 67, 1, 6, 78, 2, 12, 138, 0, 8, 138, 1, 16, 
/* out0167_had-eta7-phi8*/	6, 66, 0, 2, 66, 1, 4, 77, 0, 4, 77, 2, 6, 78, 1, 3, 78, 2, 1, 
/* out0168_had-eta8-phi8*/	3, 77, 0, 1, 77, 1, 7, 77, 2, 8, 
/* out0169_had-eta9-phi8*/	3, 76, 0, 11, 76, 2, 1, 77, 1, 2, 
/* out0170_had-eta10-phi8*/	2, 76, 0, 2, 76, 1, 9, 
/* out0171_had-eta11-phi8*/	5, 15, 0, 13, 15, 1, 2, 20, 8, 14, 20, 11, 2, 76, 1, 2, 
/* out0172_had-eta12-phi8*/	6, 15, 1, 14, 15, 7, 8, 19, 3, 1, 19, 9, 1, 20, 5, 1, 20, 11, 7, 
/* out0173_had-eta13-phi8*/	6, 15, 4, 1, 15, 7, 3, 19, 3, 1, 19, 8, 4, 19, 9, 15, 19, 10, 3, 
/* out0174_had-eta14-phi8*/	4, 19, 6, 2, 19, 8, 3, 19, 10, 10, 19, 11, 7, 
/* out0175_had-eta15-phi8*/	4, 18, 3, 2, 19, 5, 13, 19, 6, 1, 19, 11, 3, 
/* out0176_had-eta16-phi8*/	3, 18, 0, 1, 18, 2, 2, 18, 3, 12, 
/* out0177_had-eta17-phi8*/	3, 18, 2, 11, 18, 6, 1, 18, 10, 2, 
/* out0178_had-eta18-phi8*/	2, 18, 6, 10, 18, 7, 1, 
/* out0179_had-eta19-phi8*/	3, 18, 4, 7, 18, 5, 1, 18, 7, 1, 
/* out0180_had-eta0-phi9*/	1, 141, 1, 6, 
/* out0181_had-eta1-phi9*/	2, 140, 3, 3, 141, 1, 10, 
/* out0182_had-eta2-phi9*/	4, 69, 0, 2, 81, 1, 2, 140, 2, 5, 140, 3, 13, 
/* out0183_had-eta3-phi9*/	8, 69, 0, 10, 69, 1, 9, 80, 0, 6, 80, 2, 7, 81, 0, 4, 81, 1, 14, 139, 3, 6, 140, 2, 11, 
/* out0184_had-eta4-phi9*/	9, 68, 0, 5, 68, 1, 2, 79, 0, 6, 79, 2, 3, 80, 0, 1, 80, 1, 9, 80, 2, 9, 139, 2, 7, 139, 3, 10, 
/* out0185_had-eta5-phi9*/	6, 78, 0, 1, 79, 0, 6, 79, 1, 13, 79, 2, 10, 138, 3, 8, 139, 2, 9, 
/* out0186_had-eta6-phi9*/	6, 78, 0, 15, 78, 1, 5, 78, 2, 3, 90, 2, 2, 138, 2, 16, 138, 3, 8, 
/* out0187_had-eta7-phi9*/	3, 77, 0, 6, 78, 1, 8, 89, 2, 6, 
/* out0188_had-eta8-phi9*/	5, 77, 0, 5, 77, 1, 6, 88, 0, 1, 88, 2, 3, 89, 2, 2, 
/* out0189_had-eta9-phi9*/	3, 76, 0, 2, 77, 1, 1, 88, 2, 11, 
/* out0190_had-eta10-phi9*/	6, 20, 3, 11, 20, 9, 9, 76, 0, 1, 76, 1, 1, 88, 1, 3, 88, 2, 1, 
/* out0191_had-eta11-phi9*/	7, 20, 2, 7, 20, 3, 2, 20, 6, 3, 20, 8, 2, 20, 9, 7, 20, 10, 15, 20, 11, 3, 
/* out0192_had-eta12-phi9*/	6, 19, 3, 2, 20, 4, 4, 20, 5, 15, 20, 6, 6, 20, 10, 1, 20, 11, 4, 
/* out0193_had-eta13-phi9*/	5, 19, 0, 6, 19, 1, 1, 19, 2, 7, 19, 3, 12, 19, 10, 1, 
/* out0194_had-eta14-phi9*/	4, 19, 2, 8, 19, 6, 11, 19, 7, 1, 19, 10, 2, 
/* out0195_had-eta15-phi9*/	4, 19, 4, 11, 19, 5, 3, 19, 6, 2, 19, 7, 2, 
/* out0196_had-eta16-phi9*/	2, 18, 0, 12, 19, 4, 2, 
/* out0197_had-eta17-phi9*/	3, 18, 0, 2, 18, 1, 9, 18, 2, 2, 
/* out0198_had-eta18-phi9*/	4, 18, 1, 2, 18, 2, 1, 18, 6, 1, 18, 7, 8, 
/* out0199_had-eta19-phi9*/	4, 4, 4, 15, 4, 5, 1, 18, 4, 4, 18, 7, 3, 
/* out0200_had-eta0-phi10*/	1, 145, 0, 6, 
/* out0201_had-eta1-phi10*/	2, 144, 0, 3, 145, 0, 10, 
/* out0202_had-eta2-phi10*/	2, 144, 0, 13, 144, 1, 5, 
/* out0203_had-eta3-phi10*/	7, 80, 0, 6, 81, 0, 12, 92, 0, 5, 92, 1, 2, 92, 2, 15, 143, 0, 6, 144, 1, 11, 
/* out0204_had-eta4-phi10*/	10, 79, 0, 1, 80, 0, 3, 80, 1, 7, 91, 0, 7, 91, 1, 1, 91, 2, 12, 92, 1, 4, 92, 2, 1, 143, 0, 10, 143, 1, 7, 
/* out0205_had-eta5-phi10*/	8, 79, 0, 3, 79, 1, 3, 90, 0, 7, 90, 2, 5, 91, 1, 7, 91, 2, 4, 142, 0, 8, 143, 1, 9, 
/* out0206_had-eta6-phi10*/	6, 89, 0, 2, 90, 0, 2, 90, 1, 11, 90, 2, 9, 142, 0, 8, 142, 1, 16, 
/* out0207_had-eta7-phi10*/	3, 89, 0, 10, 89, 1, 3, 89, 2, 7, 
/* out0208_had-eta8-phi10*/	3, 88, 0, 6, 89, 1, 9, 89, 2, 1, 
/* out0209_had-eta9-phi10*/	3, 88, 0, 7, 88, 1, 5, 88, 2, 1, 
/* out0210_had-eta10-phi10*/	4, 20, 0, 11, 20, 3, 2, 28, 2, 2, 88, 1, 7, 
/* out0211_had-eta11-phi10*/	6, 20, 0, 5, 20, 1, 14, 20, 2, 9, 20, 3, 1, 20, 6, 4, 20, 7, 3, 
/* out0212_had-eta12-phi10*/	5, 7, 8, 5, 7, 9, 1, 20, 4, 11, 20, 6, 3, 20, 7, 11, 
/* out0213_had-eta13-phi10*/	5, 7, 8, 9, 7, 11, 2, 19, 0, 10, 19, 1, 3, 20, 4, 1, 
/* out0214_had-eta14-phi10*/	4, 7, 11, 1, 19, 1, 12, 19, 2, 1, 19, 7, 8, 
/* out0215_had-eta15-phi10*/	4, 6, 8, 3, 6, 9, 6, 19, 4, 3, 19, 7, 5, 
/* out0216_had-eta16-phi10*/	3, 6, 8, 12, 6, 9, 1, 6, 11, 2, 
/* out0217_had-eta17-phi10*/	4, 6, 8, 1, 6, 11, 8, 18, 0, 1, 18, 1, 3, 
/* out0218_had-eta18-phi10*/	6, 4, 3, 1, 4, 5, 3, 6, 5, 1, 6, 11, 1, 18, 1, 2, 18, 7, 3, 
/* out0219_had-eta19-phi10*/	2, 4, 4, 1, 4, 5, 10, 
/* out0220_had-eta0-phi11*/	1, 145, 1, 6, 
/* out0221_had-eta1-phi11*/	2, 144, 3, 3, 145, 1, 10, 
/* out0222_had-eta2-phi11*/	2, 144, 2, 5, 144, 3, 13, 
/* out0223_had-eta3-phi11*/	4, 92, 0, 11, 92, 1, 6, 143, 3, 6, 144, 2, 11, 
/* out0224_had-eta4-phi11*/	6, 31, 0, 1, 91, 0, 9, 91, 1, 2, 92, 1, 4, 143, 2, 7, 143, 3, 10, 
/* out0225_had-eta5-phi11*/	7, 31, 0, 3, 31, 1, 1, 31, 2, 15, 90, 0, 4, 91, 1, 6, 142, 3, 8, 143, 2, 9, 
/* out0226_had-eta6-phi11*/	8, 30, 0, 4, 30, 2, 8, 31, 1, 2, 31, 2, 1, 90, 0, 3, 90, 1, 5, 142, 2, 16, 142, 3, 8, 
/* out0227_had-eta7-phi11*/	5, 29, 0, 2, 30, 1, 4, 30, 2, 8, 89, 0, 4, 89, 1, 2, 
/* out0228_had-eta8-phi11*/	3, 29, 0, 2, 29, 2, 12, 89, 1, 2, 
/* out0229_had-eta9-phi11*/	6, 28, 0, 2, 28, 2, 1, 29, 1, 4, 29, 2, 4, 88, 0, 2, 88, 1, 1, 
/* out0230_had-eta10-phi11*/	2, 28, 0, 2, 28, 2, 9, 
/* out0231_had-eta11-phi11*/	5, 7, 3, 3, 20, 1, 2, 20, 7, 1, 28, 1, 4, 28, 2, 4, 
/* out0232_had-eta12-phi11*/	5, 7, 2, 3, 7, 3, 9, 7, 9, 14, 7, 10, 4, 20, 7, 1, 
/* out0233_had-eta13-phi11*/	6, 7, 5, 1, 7, 6, 4, 7, 8, 2, 7, 9, 1, 7, 10, 12, 7, 11, 8, 
/* out0234_had-eta14-phi11*/	4, 6, 3, 5, 6, 9, 1, 7, 5, 11, 7, 11, 5, 
/* out0235_had-eta15-phi11*/	4, 6, 2, 3, 6, 3, 6, 6, 9, 7, 6, 10, 3, 
/* out0236_had-eta16-phi11*/	5, 6, 2, 1, 6, 6, 1, 6, 9, 1, 6, 10, 12, 6, 11, 1, 
/* out0237_had-eta17-phi11*/	4, 6, 5, 6, 6, 6, 3, 6, 10, 1, 6, 11, 4, 
/* out0238_had-eta18-phi11*/	2, 4, 3, 6, 6, 5, 5, 
/* out0239_had-eta19-phi11*/	4, 4, 2, 4, 4, 3, 5, 4, 5, 2, 4, 6, 16, 
/* out0240_had-eta0-phi12*/	1, 149, 0, 6, 
/* out0241_had-eta1-phi12*/	2, 148, 0, 3, 149, 0, 10, 
/* out0242_had-eta2-phi12*/	2, 148, 0, 13, 148, 1, 5, 
/* out0243_had-eta3-phi12*/	4, 41, 0, 4, 41, 2, 14, 147, 0, 6, 148, 1, 11, 
/* out0244_had-eta4-phi12*/	7, 31, 0, 1, 40, 0, 2, 40, 2, 10, 41, 1, 2, 41, 2, 2, 147, 0, 10, 147, 1, 7, 
/* out0245_had-eta5-phi12*/	8, 31, 0, 11, 31, 1, 9, 39, 0, 1, 39, 2, 3, 40, 1, 1, 40, 2, 5, 146, 0, 8, 147, 1, 9, 
/* out0246_had-eta6-phi12*/	5, 30, 0, 12, 31, 1, 4, 39, 2, 8, 146, 0, 8, 146, 1, 16, 
/* out0247_had-eta7-phi12*/	3, 29, 0, 2, 30, 1, 12, 38, 2, 6, 
/* out0248_had-eta8-phi12*/	3, 29, 0, 10, 29, 1, 5, 38, 2, 1, 
/* out0249_had-eta9-phi12*/	3, 28, 0, 3, 29, 1, 7, 37, 2, 3, 
/* out0250_had-eta10-phi12*/	2, 28, 0, 8, 28, 1, 3, 
/* out0251_had-eta11-phi12*/	3, 7, 0, 3, 13, 8, 3, 28, 1, 8, 
/* out0252_had-eta12-phi12*/	5, 7, 0, 12, 7, 1, 7, 7, 2, 8, 7, 3, 4, 13, 8, 1, 
/* out0253_had-eta13-phi12*/	6, 7, 1, 1, 7, 2, 5, 7, 4, 1, 7, 5, 1, 7, 6, 12, 7, 7, 7, 
/* out0254_had-eta14-phi12*/	4, 6, 0, 6, 6, 3, 1, 7, 4, 12, 7, 5, 3, 
/* out0255_had-eta15-phi12*/	4, 6, 0, 6, 6, 1, 3, 6, 2, 6, 6, 3, 4, 
/* out0256_had-eta16-phi12*/	2, 6, 2, 6, 6, 6, 8, 
/* out0257_had-eta17-phi12*/	4, 6, 4, 4, 6, 5, 3, 6, 6, 4, 6, 7, 1, 
/* out0258_had-eta18-phi12*/	4, 4, 0, 5, 4, 3, 1, 6, 4, 4, 6, 5, 1, 
/* out0259_had-eta19-phi12*/	4, 4, 0, 3, 4, 1, 1, 4, 2, 5, 4, 3, 3, 
/* out0260_had-eta0-phi13*/	1, 149, 1, 6, 
/* out0261_had-eta1-phi13*/	2, 148, 3, 3, 149, 1, 10, 
/* out0262_had-eta2-phi13*/	2, 148, 2, 5, 148, 3, 13, 
/* out0263_had-eta3-phi13*/	8, 41, 0, 12, 41, 1, 9, 52, 0, 2, 52, 2, 4, 53, 0, 4, 53, 1, 16, 147, 3, 6, 148, 2, 11, 
/* out0264_had-eta4-phi13*/	8, 40, 0, 14, 40, 1, 4, 40, 2, 1, 41, 1, 5, 51, 2, 1, 52, 2, 10, 147, 2, 7, 147, 3, 10, 
/* out0265_had-eta5-phi13*/	6, 39, 0, 12, 39, 2, 1, 40, 1, 11, 51, 2, 6, 146, 3, 8, 147, 2, 9, 
/* out0266_had-eta6-phi13*/	7, 38, 0, 2, 39, 0, 3, 39, 1, 15, 39, 2, 4, 50, 2, 1, 146, 2, 16, 146, 3, 8, 
/* out0267_had-eta7-phi13*/	3, 38, 0, 11, 38, 1, 3, 38, 2, 6, 
/* out0268_had-eta8-phi13*/	4, 37, 0, 5, 37, 2, 1, 38, 1, 8, 38, 2, 3, 
/* out0269_had-eta9-phi13*/	3, 37, 0, 3, 37, 1, 2, 37, 2, 9, 
/* out0270_had-eta10-phi13*/	6, 13, 3, 10, 13, 9, 3, 28, 0, 1, 28, 1, 1, 37, 1, 4, 37, 2, 3, 
/* out0271_had-eta11-phi13*/	6, 13, 2, 2, 13, 3, 2, 13, 8, 8, 13, 9, 13, 13, 10, 11, 13, 11, 1, 
/* out0272_had-eta12-phi13*/	6, 7, 0, 1, 7, 1, 6, 13, 5, 4, 13, 8, 4, 13, 10, 3, 13, 11, 15, 
/* out0273_had-eta13-phi13*/	5, 7, 1, 2, 7, 4, 1, 7, 7, 9, 11, 3, 2, 11, 9, 11, 
/* out0274_had-eta14-phi13*/	6, 6, 0, 1, 7, 4, 2, 11, 8, 14, 11, 9, 4, 11, 10, 1, 11, 11, 2, 
/* out0275_had-eta15-phi13*/	4, 6, 0, 3, 6, 1, 7, 11, 8, 2, 11, 11, 6, 
/* out0276_had-eta16-phi13*/	2, 6, 1, 5, 6, 7, 10, 
/* out0277_had-eta17-phi13*/	4, 5, 8, 3, 5, 9, 1, 6, 4, 6, 6, 7, 4, 
/* out0278_had-eta18-phi13*/	3, 4, 0, 3, 5, 8, 6, 6, 4, 2, 
/* out0279_had-eta19-phi13*/	3, 4, 0, 5, 4, 1, 7, 4, 2, 7, 
/* out0280_had-eta0-phi14*/	1, 153, 0, 6, 
/* out0281_had-eta1-phi14*/	2, 152, 0, 3, 153, 0, 10, 
/* out0282_had-eta2-phi14*/	4, 53, 0, 1, 63, 0, 2, 152, 0, 13, 152, 1, 5, 
/* out0283_had-eta3-phi14*/	7, 52, 0, 13, 53, 0, 11, 63, 0, 2, 63, 1, 1, 63, 2, 16, 151, 0, 6, 152, 1, 11, 
/* out0284_had-eta4-phi14*/	7, 51, 0, 9, 52, 0, 1, 52, 1, 16, 52, 2, 2, 62, 2, 7, 151, 0, 10, 151, 1, 7, 
/* out0285_had-eta5-phi14*/	6, 50, 0, 1, 51, 0, 6, 51, 1, 14, 51, 2, 9, 150, 0, 8, 151, 1, 9, 
/* out0286_had-eta6-phi14*/	6, 39, 1, 1, 50, 0, 9, 50, 1, 2, 50, 2, 11, 150, 0, 8, 150, 1, 16, 
/* out0287_had-eta7-phi14*/	6, 38, 0, 3, 38, 1, 3, 49, 0, 3, 49, 2, 2, 50, 1, 4, 50, 2, 4, 
/* out0288_had-eta8-phi14*/	3, 37, 0, 3, 38, 1, 2, 49, 2, 11, 
/* out0289_had-eta9-phi14*/	4, 37, 0, 5, 37, 1, 6, 48, 2, 1, 49, 2, 1, 
/* out0290_had-eta10-phi14*/	5, 13, 0, 16, 13, 1, 1, 13, 3, 3, 37, 1, 4, 48, 2, 3, 
/* out0291_had-eta11-phi14*/	6, 13, 1, 8, 13, 2, 14, 13, 3, 1, 13, 6, 9, 13, 7, 3, 13, 10, 2, 
/* out0292_had-eta12-phi14*/	5, 11, 0, 2, 13, 4, 9, 13, 5, 12, 13, 6, 7, 13, 7, 2, 
/* out0293_had-eta13-phi14*/	5, 11, 0, 4, 11, 2, 7, 11, 3, 14, 11, 9, 1, 11, 10, 1, 
/* out0294_had-eta14-phi14*/	4, 11, 2, 3, 11, 6, 4, 11, 10, 13, 11, 11, 1, 
/* out0295_had-eta15-phi14*/	4, 11, 5, 9, 11, 6, 2, 11, 10, 1, 11, 11, 7, 
/* out0296_had-eta16-phi14*/	5, 5, 3, 7, 5, 9, 6, 6, 1, 1, 6, 7, 1, 11, 5, 2, 
/* out0297_had-eta17-phi14*/	3, 5, 8, 1, 5, 9, 9, 5, 10, 3, 
/* out0298_had-eta18-phi14*/	3, 5, 8, 5, 5, 10, 2, 5, 11, 4, 
/* out0299_had-eta19-phi14*/	3, 4, 1, 8, 5, 8, 1, 5, 11, 6, 
/* out0300_had-eta0-phi15*/	1, 153, 1, 6, 
/* out0301_had-eta1-phi15*/	2, 152, 3, 3, 153, 1, 10, 
/* out0302_had-eta2-phi15*/	3, 63, 0, 4, 152, 2, 5, 152, 3, 13, 
/* out0303_had-eta3-phi15*/	7, 62, 0, 5, 63, 0, 8, 63, 1, 15, 106, 0, 3, 106, 2, 11, 151, 3, 6, 152, 2, 11, 
/* out0304_had-eta4-phi15*/	5, 62, 0, 11, 62, 1, 14, 62, 2, 9, 151, 2, 7, 151, 3, 10, 
/* out0305_had-eta5-phi15*/	8, 51, 0, 1, 51, 1, 2, 61, 0, 10, 61, 1, 2, 61, 2, 13, 62, 1, 1, 150, 3, 8, 151, 2, 9, 
/* out0306_had-eta6-phi15*/	8, 50, 0, 6, 50, 1, 6, 60, 0, 2, 60, 2, 4, 61, 1, 3, 61, 2, 3, 150, 2, 16, 150, 3, 8, 
/* out0307_had-eta7-phi15*/	3, 49, 0, 10, 50, 1, 4, 60, 2, 6, 
/* out0308_had-eta8-phi15*/	3, 49, 0, 3, 49, 1, 12, 49, 2, 2, 
/* out0309_had-eta9-phi15*/	3, 48, 0, 9, 48, 2, 3, 49, 1, 2, 
/* out0310_had-eta10-phi15*/	2, 48, 1, 3, 48, 2, 8, 
/* out0311_had-eta11-phi15*/	6, 12, 3, 5, 12, 9, 9, 13, 1, 7, 13, 7, 10, 48, 1, 1, 48, 2, 1, 
/* out0312_had-eta12-phi15*/	6, 11, 0, 2, 12, 8, 14, 12, 9, 6, 12, 11, 1, 13, 4, 7, 13, 7, 1, 
/* out0313_had-eta13-phi15*/	5, 11, 0, 8, 11, 1, 12, 11, 2, 3, 12, 8, 2, 12, 11, 2, 
/* out0314_had-eta14-phi15*/	5, 11, 1, 1, 11, 2, 3, 11, 4, 1, 11, 6, 9, 11, 7, 8, 
/* out0315_had-eta15-phi15*/	4, 5, 0, 2, 11, 4, 11, 11, 5, 5, 11, 6, 1, 
/* out0316_had-eta16-phi15*/	3, 5, 0, 5, 5, 2, 2, 5, 3, 9, 
/* out0317_had-eta17-phi15*/	2, 5, 2, 7, 5, 10, 5, 
/* out0318_had-eta18-phi15*/	4, 5, 5, 2, 5, 6, 4, 5, 10, 6, 5, 11, 1, 
/* out0319_had-eta19-phi15*/	2, 5, 5, 5, 5, 11, 5, 
/* out0320_had-eta0-phi16*/	1, 157, 0, 6, 
/* out0321_had-eta1-phi16*/	2, 156, 0, 3, 157, 0, 10, 
/* out0322_had-eta2-phi16*/	4, 107, 0, 2, 107, 1, 11, 156, 0, 13, 156, 1, 5, 
/* out0323_had-eta3-phi16*/	9, 105, 0, 1, 105, 2, 5, 106, 0, 13, 106, 1, 14, 106, 2, 4, 107, 0, 3, 107, 1, 5, 155, 0, 6, 156, 1, 11, 
/* out0324_had-eta4-phi16*/	9, 62, 1, 1, 104, 0, 14, 104, 1, 5, 104, 2, 13, 105, 2, 1, 106, 1, 2, 106, 2, 1, 155, 0, 10, 155, 1, 7, 
/* out0325_had-eta5-phi16*/	8, 61, 0, 6, 61, 1, 8, 103, 0, 3, 103, 2, 6, 104, 1, 4, 104, 2, 3, 154, 0, 8, 155, 1, 9, 
/* out0326_had-eta6-phi16*/	7, 60, 0, 14, 60, 1, 2, 60, 2, 1, 61, 1, 3, 103, 2, 5, 154, 0, 8, 154, 1, 16, 
/* out0327_had-eta7-phi16*/	3, 59, 0, 3, 60, 1, 11, 60, 2, 5, 
/* out0328_had-eta8-phi16*/	3, 49, 1, 2, 59, 0, 3, 59, 2, 11, 
/* out0329_had-eta9-phi16*/	3, 48, 0, 7, 48, 1, 2, 59, 2, 5, 
/* out0330_had-eta10-phi16*/	3, 12, 0, 1, 48, 1, 10, 70, 2, 1, 
/* out0331_had-eta11-phi16*/	6, 12, 0, 12, 12, 1, 1, 12, 2, 10, 12, 3, 11, 12, 9, 1, 12, 10, 1, 
/* out0332_had-eta12-phi16*/	5, 12, 2, 4, 12, 5, 1, 12, 6, 9, 12, 10, 15, 12, 11, 4, 
/* out0333_had-eta13-phi16*/	6, 11, 1, 3, 11, 7, 1, 12, 5, 9, 12, 11, 9, 16, 3, 3, 16, 9, 1, 
/* out0334_had-eta14-phi16*/	4, 11, 4, 1, 11, 7, 7, 16, 8, 1, 16, 9, 10, 
/* out0335_had-eta15-phi16*/	3, 5, 0, 2, 11, 4, 3, 16, 8, 11, 
/* out0336_had-eta16-phi16*/	4, 5, 0, 7, 5, 1, 6, 5, 2, 1, 16, 8, 1, 
/* out0337_had-eta17-phi16*/	4, 5, 1, 2, 5, 2, 6, 5, 6, 5, 5, 7, 1, 
/* out0338_had-eta18-phi16*/	4, 5, 4, 1, 5, 5, 2, 5, 6, 7, 5, 7, 1, 
/* out0339_had-eta19-phi16*/	2, 5, 4, 3, 5, 5, 7, 
/* out0340_had-eta0-phi17*/	1, 157, 1, 6, 
/* out0341_had-eta1-phi17*/	2, 156, 3, 3, 157, 1, 10, 
/* out0342_had-eta2-phi17*/	3, 107, 0, 7, 156, 2, 5, 156, 3, 13, 
/* out0343_had-eta3-phi17*/	6, 105, 0, 15, 105, 1, 10, 105, 2, 7, 107, 0, 4, 155, 3, 6, 156, 2, 11, 
/* out0344_had-eta4-phi17*/	8, 104, 0, 2, 104, 1, 6, 105, 1, 6, 105, 2, 3, 119, 0, 8, 119, 2, 11, 155, 2, 7, 155, 3, 10, 
/* out0345_had-eta5-phi17*/	7, 103, 0, 13, 103, 1, 7, 103, 2, 2, 104, 1, 1, 119, 2, 5, 154, 3, 8, 155, 2, 9, 
/* out0346_had-eta6-phi17*/	7, 60, 1, 1, 103, 1, 9, 103, 2, 3, 115, 0, 7, 115, 2, 2, 154, 2, 16, 154, 3, 8, 
/* out0347_had-eta7-phi17*/	3, 59, 0, 4, 60, 1, 2, 115, 2, 13, 
/* out0348_had-eta8-phi17*/	2, 59, 0, 6, 59, 1, 10, 
/* out0349_had-eta9-phi17*/	3, 59, 1, 6, 70, 0, 7, 70, 2, 1, 
/* out0350_had-eta10-phi17*/	2, 70, 0, 1, 70, 2, 11, 
/* out0351_had-eta11-phi17*/	5, 12, 0, 3, 12, 1, 15, 12, 2, 2, 12, 7, 5, 70, 2, 3, 
/* out0352_had-eta12-phi17*/	4, 12, 4, 10, 12, 5, 2, 12, 6, 7, 12, 7, 11, 
/* out0353_had-eta13-phi17*/	4, 12, 4, 6, 12, 5, 4, 16, 0, 7, 16, 3, 9, 
/* out0354_had-eta14-phi17*/	4, 16, 2, 7, 16, 3, 4, 16, 9, 4, 16, 10, 7, 
/* out0355_had-eta15-phi17*/	4, 16, 8, 2, 16, 9, 1, 16, 10, 8, 16, 11, 7, 
/* out0356_had-eta16-phi17*/	3, 5, 1, 6, 16, 8, 1, 16, 11, 8, 
/* out0357_had-eta17-phi17*/	2, 5, 1, 2, 5, 7, 11, 
/* out0358_had-eta18-phi17*/	2, 5, 4, 7, 5, 7, 3, 
/* out0359_had-eta19-phi17*/	1, 5, 4, 5, 
/* out0360_had-eta0-phi18*/	1, 161, 0, 6, 
/* out0361_had-eta1-phi18*/	2, 160, 0, 3, 161, 0, 10, 
/* out0362_had-eta2-phi18*/	3, 121, 1, 7, 160, 0, 13, 160, 1, 5, 
/* out0363_had-eta3-phi18*/	6, 120, 0, 15, 120, 1, 7, 120, 2, 10, 121, 1, 4, 159, 0, 6, 160, 1, 11, 
/* out0364_had-eta4-phi18*/	8, 117, 0, 2, 117, 2, 6, 119, 0, 8, 119, 1, 10, 120, 1, 3, 120, 2, 6, 159, 0, 10, 159, 1, 7, 
/* out0365_had-eta5-phi18*/	7, 116, 0, 13, 116, 1, 2, 116, 2, 7, 117, 2, 1, 119, 1, 6, 158, 0, 8, 159, 1, 9, 
/* out0366_had-eta6-phi18*/	7, 72, 2, 1, 115, 0, 8, 115, 1, 2, 116, 1, 3, 116, 2, 9, 158, 0, 8, 158, 1, 16, 
/* out0367_had-eta7-phi18*/	5, 71, 0, 4, 72, 2, 2, 115, 0, 1, 115, 1, 14, 115, 2, 1, 
/* out0368_had-eta8-phi18*/	2, 71, 0, 6, 71, 2, 10, 
/* out0369_had-eta9-phi18*/	3, 70, 0, 7, 70, 1, 1, 71, 2, 6, 
/* out0370_had-eta10-phi18*/	2, 70, 0, 1, 70, 1, 10, 
/* out0371_had-eta11-phi18*/	5, 17, 0, 3, 17, 2, 2, 17, 3, 15, 17, 9, 5, 70, 1, 3, 
/* out0372_had-eta12-phi18*/	4, 17, 8, 10, 17, 9, 11, 17, 10, 7, 17, 11, 2, 
/* out0373_had-eta13-phi18*/	4, 16, 0, 9, 16, 1, 8, 17, 8, 6, 17, 11, 4, 
/* out0374_had-eta14-phi18*/	4, 16, 1, 4, 16, 2, 9, 16, 6, 7, 16, 7, 2, 
/* out0375_had-eta15-phi18*/	5, 16, 4, 1, 16, 5, 7, 16, 6, 9, 16, 7, 1, 16, 10, 1, 
/* out0376_had-eta16-phi18*/	3, 16, 5, 9, 16, 11, 1, 21, 3, 6, 
/* out0377_had-eta17-phi18*/	2, 21, 3, 2, 21, 9, 11, 
/* out0378_had-eta18-phi18*/	2, 21, 8, 7, 21, 9, 3, 
/* out0379_had-eta19-phi18*/	1, 21, 8, 5, 
/* out0380_had-eta0-phi19*/	1, 161, 1, 6, 
/* out0381_had-eta1-phi19*/	2, 160, 3, 3, 161, 1, 10, 
/* out0382_had-eta2-phi19*/	4, 121, 0, 11, 121, 1, 2, 160, 2, 5, 160, 3, 13, 
/* out0383_had-eta3-phi19*/	9, 118, 0, 13, 118, 1, 4, 118, 2, 14, 120, 0, 1, 120, 1, 5, 121, 0, 5, 121, 1, 3, 159, 3, 6, 160, 2, 11, 
/* out0384_had-eta4-phi19*/	9, 74, 2, 1, 117, 0, 14, 117, 1, 13, 117, 2, 5, 118, 1, 1, 118, 2, 2, 120, 1, 1, 159, 2, 7, 159, 3, 10, 
/* out0385_had-eta5-phi19*/	8, 73, 0, 6, 73, 2, 8, 116, 0, 3, 116, 1, 6, 117, 1, 3, 117, 2, 4, 158, 3, 8, 159, 2, 9, 
/* out0386_had-eta6-phi19*/	7, 72, 0, 14, 72, 1, 1, 72, 2, 2, 73, 2, 3, 116, 1, 5, 158, 2, 16, 158, 3, 8, 
/* out0387_had-eta7-phi19*/	3, 71, 0, 3, 72, 1, 5, 72, 2, 11, 
/* out0388_had-eta8-phi19*/	3, 71, 0, 3, 71, 1, 11, 83, 2, 2, 
/* out0389_had-eta9-phi19*/	3, 71, 1, 5, 82, 0, 7, 82, 2, 2, 
/* out0390_had-eta10-phi19*/	3, 17, 0, 1, 70, 1, 2, 82, 2, 10, 
/* out0391_had-eta11-phi19*/	6, 17, 0, 12, 17, 1, 11, 17, 2, 10, 17, 3, 1, 17, 6, 1, 17, 7, 1, 
/* out0392_had-eta12-phi19*/	5, 17, 2, 4, 17, 5, 4, 17, 6, 15, 17, 10, 9, 17, 11, 1, 
/* out0393_had-eta13-phi19*/	6, 16, 1, 3, 16, 7, 1, 17, 5, 9, 17, 11, 9, 22, 3, 3, 22, 9, 1, 
/* out0394_had-eta14-phi19*/	5, 16, 1, 1, 16, 4, 1, 16, 7, 12, 22, 8, 1, 22, 9, 7, 
/* out0395_had-eta15-phi19*/	3, 16, 4, 13, 21, 0, 2, 22, 8, 3, 
/* out0396_had-eta16-phi19*/	4, 16, 4, 1, 21, 0, 7, 21, 2, 1, 21, 3, 6, 
/* out0397_had-eta17-phi19*/	4, 21, 2, 6, 21, 3, 2, 21, 9, 1, 21, 10, 5, 
/* out0398_had-eta18-phi19*/	4, 21, 8, 1, 21, 9, 1, 21, 10, 7, 21, 11, 2, 
/* out0399_had-eta19-phi19*/	2, 21, 8, 3, 21, 11, 7, 
/* out0400_had-eta0-phi20*/	1, 165, 0, 6, 
/* out0401_had-eta1-phi20*/	2, 164, 0, 3, 165, 0, 10, 
/* out0402_had-eta2-phi20*/	3, 75, 0, 4, 164, 0, 13, 164, 1, 5, 
/* out0403_had-eta3-phi20*/	7, 74, 0, 5, 75, 0, 8, 75, 2, 15, 118, 0, 3, 118, 1, 11, 163, 0, 6, 164, 1, 11, 
/* out0404_had-eta4-phi20*/	5, 74, 0, 11, 74, 1, 9, 74, 2, 14, 163, 0, 10, 163, 1, 7, 
/* out0405_had-eta5-phi20*/	8, 73, 0, 10, 73, 1, 13, 73, 2, 2, 74, 2, 1, 85, 0, 1, 85, 2, 2, 162, 0, 8, 163, 1, 9, 
/* out0406_had-eta6-phi20*/	8, 72, 0, 2, 72, 1, 4, 73, 1, 3, 73, 2, 3, 84, 0, 6, 84, 2, 6, 162, 0, 8, 162, 1, 16, 
/* out0407_had-eta7-phi20*/	3, 72, 1, 6, 83, 0, 10, 84, 2, 4, 
/* out0408_had-eta8-phi20*/	3, 83, 0, 3, 83, 1, 2, 83, 2, 12, 
/* out0409_had-eta9-phi20*/	3, 82, 0, 9, 82, 1, 3, 83, 2, 2, 
/* out0410_had-eta10-phi20*/	2, 82, 1, 8, 82, 2, 3, 
/* out0411_had-eta11-phi20*/	6, 17, 1, 5, 17, 7, 9, 23, 3, 7, 23, 9, 10, 82, 1, 1, 82, 2, 1, 
/* out0412_had-eta12-phi20*/	6, 17, 4, 14, 17, 5, 1, 17, 7, 6, 22, 0, 2, 23, 8, 7, 23, 9, 1, 
/* out0413_had-eta13-phi20*/	5, 17, 4, 2, 17, 5, 2, 22, 0, 8, 22, 2, 3, 22, 3, 12, 
/* out0414_had-eta14-phi20*/	5, 22, 2, 3, 22, 3, 1, 22, 8, 1, 22, 9, 8, 22, 10, 9, 
/* out0415_had-eta15-phi20*/	4, 21, 0, 2, 22, 8, 11, 22, 10, 1, 22, 11, 5, 
/* out0416_had-eta16-phi20*/	3, 21, 0, 5, 21, 1, 9, 21, 2, 2, 
/* out0417_had-eta17-phi20*/	2, 21, 2, 7, 21, 6, 5, 
/* out0418_had-eta18-phi20*/	4, 21, 5, 1, 21, 6, 6, 21, 10, 4, 21, 11, 2, 
/* out0419_had-eta19-phi20*/	2, 21, 5, 5, 21, 11, 5, 
/* out0420_had-eta0-phi21*/	1, 165, 1, 6, 
/* out0421_had-eta1-phi21*/	2, 164, 3, 3, 165, 1, 10, 
/* out0422_had-eta2-phi21*/	4, 75, 0, 2, 87, 1, 1, 164, 2, 5, 164, 3, 13, 
/* out0423_had-eta3-phi21*/	7, 75, 0, 2, 75, 1, 16, 75, 2, 1, 86, 0, 13, 87, 1, 11, 163, 3, 6, 164, 2, 11, 
/* out0424_had-eta4-phi21*/	7, 74, 1, 7, 85, 0, 9, 86, 0, 1, 86, 1, 2, 86, 2, 16, 163, 2, 7, 163, 3, 10, 
/* out0425_had-eta5-phi21*/	6, 84, 0, 1, 85, 0, 6, 85, 1, 9, 85, 2, 14, 162, 3, 8, 163, 2, 9, 
/* out0426_had-eta6-phi21*/	6, 84, 0, 9, 84, 1, 11, 84, 2, 2, 95, 2, 1, 162, 2, 16, 162, 3, 8, 
/* out0427_had-eta7-phi21*/	6, 83, 0, 3, 83, 1, 2, 84, 1, 4, 84, 2, 4, 94, 0, 3, 94, 2, 3, 
/* out0428_had-eta8-phi21*/	3, 83, 1, 11, 93, 0, 3, 94, 2, 2, 
/* out0429_had-eta9-phi21*/	4, 82, 1, 1, 83, 1, 1, 93, 0, 5, 93, 2, 6, 
/* out0430_had-eta10-phi21*/	5, 23, 0, 16, 23, 1, 3, 23, 3, 1, 82, 1, 3, 93, 2, 4, 
/* out0431_had-eta11-phi21*/	6, 23, 1, 1, 23, 2, 14, 23, 3, 8, 23, 6, 2, 23, 9, 3, 23, 10, 9, 
/* out0432_had-eta12-phi21*/	5, 22, 0, 2, 23, 8, 9, 23, 9, 2, 23, 10, 7, 23, 11, 12, 
/* out0433_had-eta13-phi21*/	5, 22, 0, 4, 22, 1, 14, 22, 2, 7, 22, 6, 1, 22, 7, 1, 
/* out0434_had-eta14-phi21*/	4, 22, 2, 3, 22, 5, 1, 22, 6, 13, 22, 10, 4, 
/* out0435_had-eta15-phi21*/	4, 22, 5, 7, 22, 6, 1, 22, 10, 2, 22, 11, 9, 
/* out0436_had-eta16-phi21*/	3, 21, 1, 7, 21, 7, 6, 22, 11, 2, 
/* out0437_had-eta17-phi21*/	3, 21, 4, 1, 21, 6, 3, 21, 7, 9, 
/* out0438_had-eta18-phi21*/	3, 21, 4, 5, 21, 5, 4, 21, 6, 2, 
/* out0439_had-eta19-phi21*/	2, 21, 4, 1, 21, 5, 6, 
/* out0440_had-eta0-phi22*/	1, 169, 0, 6, 
/* out0441_had-eta1-phi22*/	2, 168, 0, 3, 169, 0, 10, 
/* out0442_had-eta2-phi22*/	2, 168, 0, 13, 168, 1, 5, 
/* out0443_had-eta3-phi22*/	8, 86, 0, 2, 86, 1, 4, 87, 0, 16, 87, 1, 4, 97, 0, 12, 97, 2, 9, 167, 0, 6, 168, 1, 11, 
/* out0444_had-eta4-phi22*/	8, 85, 1, 1, 86, 1, 10, 96, 0, 14, 96, 1, 1, 96, 2, 4, 97, 2, 5, 167, 0, 10, 167, 1, 7, 
/* out0445_had-eta5-phi22*/	6, 85, 1, 6, 95, 0, 12, 95, 1, 1, 96, 2, 11, 166, 0, 8, 167, 1, 9, 
/* out0446_had-eta6-phi22*/	7, 84, 1, 1, 94, 0, 2, 95, 0, 3, 95, 1, 4, 95, 2, 15, 166, 0, 8, 166, 1, 16, 
/* out0447_had-eta7-phi22*/	3, 94, 0, 11, 94, 1, 6, 94, 2, 3, 
/* out0448_had-eta8-phi22*/	4, 93, 0, 5, 93, 1, 1, 94, 1, 3, 94, 2, 8, 
/* out0449_had-eta9-phi22*/	3, 93, 0, 3, 93, 1, 9, 93, 2, 2, 
/* out0450_had-eta10-phi22*/	4, 23, 1, 10, 23, 7, 3, 93, 1, 3, 93, 2, 4, 
/* out0451_had-eta11-phi22*/	6, 23, 1, 2, 23, 2, 2, 23, 4, 8, 23, 5, 1, 23, 6, 11, 23, 7, 13, 
/* out0452_had-eta12-phi22*/	4, 23, 4, 4, 23, 5, 15, 23, 6, 3, 23, 11, 4, 
/* out0453_had-eta13-phi22*/	2, 22, 1, 2, 22, 7, 11, 
/* out0454_had-eta14-phi22*/	4, 22, 4, 14, 22, 5, 2, 22, 6, 1, 22, 7, 4, 
/* out0455_had-eta15-phi22*/	2, 22, 4, 2, 22, 5, 6, 
/* out0456_had-eta16-phi22*/	0, 
/* out0457_had-eta17-phi22*/	2, 21, 4, 3, 21, 7, 1, 
/* out0458_had-eta18-phi22*/	1, 21, 4, 6, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	1, 169, 1, 6, 
/* out0461_had-eta1-phi23*/	2, 168, 3, 3, 169, 1, 10, 
/* out0462_had-eta2-phi23*/	2, 168, 2, 5, 168, 3, 13, 
/* out0463_had-eta3-phi23*/	4, 97, 0, 4, 97, 1, 14, 167, 3, 6, 168, 2, 11, 
/* out0464_had-eta4-phi23*/	6, 96, 0, 2, 96, 1, 10, 97, 1, 2, 97, 2, 2, 167, 2, 7, 167, 3, 10, 
/* out0465_had-eta5-phi23*/	6, 95, 0, 1, 95, 1, 3, 96, 1, 5, 96, 2, 1, 166, 3, 8, 167, 2, 9, 
/* out0466_had-eta6-phi23*/	3, 95, 1, 8, 166, 2, 16, 166, 3, 8, 
/* out0467_had-eta7-phi23*/	1, 94, 1, 6, 
/* out0468_had-eta8-phi23*/	1, 94, 1, 1, 
/* out0469_had-eta9-phi23*/	1, 93, 1, 3, 
/* out0470_had-eta10-phi23*/	0, 
/* out0471_had-eta11-phi23*/	1, 23, 4, 3, 
/* out0472_had-eta12-phi23*/	1, 23, 4, 1, 
/* out0473_had-eta13-phi23*/	0, 
/* out0474_had-eta14-phi23*/	0, 
/* out0475_had-eta15-phi23*/	0, 
/* out0476_had-eta16-phi23*/	0, 
/* out0477_had-eta17-phi23*/	0, 
/* out0478_had-eta18-phi23*/	0, 
/* out0479_had-eta19-phi23*/	0, 
};