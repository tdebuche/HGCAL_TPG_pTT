parameter integer matrixH [0:6308] = {
/* num inputs = 182(in0-in181) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 10 */
//* total number of input in adders 1942 */

/* out0000_em-eta0-phi0*/	1,137,0,16,
/* out0001_em-eta1-phi0*/	1,137,1,15,
/* out0002_em-eta2-phi0*/	3,136,0,16,136,1,1,137,1,1,
/* out0003_em-eta3-phi0*/	6,59,0,4,59,1,2,60,1,2,60,2,12,135,0,2,136,1,15,
/* out0004_em-eta4-phi0*/	8,51,0,16,51,1,16,51,2,4,58,0,1,59,0,10,59,2,1,135,0,14,135,1,4,
/* out0005_em-eta5-phi0*/	5,50,1,7,51,2,12,58,0,10,134,0,5,135,1,12,
/* out0006_em-eta6-phi0*/	7,50,0,16,50,1,9,50,2,15,57,0,4,58,0,1,134,0,11,134,1,6,
/* out0007_em-eta7-phi0*/	7,49,0,1,49,1,15,49,2,1,50,2,1,57,0,4,134,1,10,134,2,7,
/* out0008_em-eta8-phi0*/	5,48,1,1,49,0,15,49,2,12,56,0,2,134,2,9,
/* out0009_em-eta9-phi0*/	4,48,0,1,48,1,14,48,2,1,56,0,1,
/* out0010_em-eta10-phi0*/	3,11,5,1,48,0,15,48,2,10,
/* out0011_em-eta11-phi0*/	8,6,2,1,6,3,11,7,2,16,7,3,16,7,4,3,10,5,2,11,5,1,48,2,1,
/* out0012_em-eta12-phi0*/	6,6,0,1,6,1,4,6,2,15,6,3,3,7,0,14,7,4,13,
/* out0013_em-eta13-phi0*/	6,3,2,1,3,3,4,6,1,7,6,4,16,7,0,2,7,1,16,
/* out0014_em-eta14-phi0*/	5,2,2,1,2,3,6,3,2,15,3,3,12,3,4,2,
/* out0015_em-eta15-phi0*/	4,2,2,12,2,3,1,3,0,12,3,4,14,
/* out0016_em-eta16-phi0*/	4,2,1,3,2,2,3,3,0,4,3,1,4,
/* out0017_em-eta17-phi0*/	4,0,4,4,1,1,1,2,4,16,3,1,11,
/* out0018_em-eta18-phi0*/	5,0,2,1,0,4,4,0,5,1,1,0,11,1,1,15,
/* out0019_em-eta19-phi0*/	6,0,0,16,0,2,4,0,3,9,1,0,3,1,3,4,1,5,4,
/* out0020_em-eta0-phi1*/	1,137,3,16,
/* out0021_em-eta1-phi1*/	1,137,2,15,
/* out0022_em-eta2-phi1*/	6,60,1,1,60,2,1,70,1,1,136,2,1,136,3,16,137,2,1,
/* out0023_em-eta3-phi1*/	7,59,1,11,60,1,13,60,2,3,70,0,14,70,1,1,135,3,2,136,2,15,
/* out0024_em-eta4-phi1*/	7,58,1,5,59,0,2,59,1,3,59,2,15,69,0,6,135,2,4,135,3,14,
/* out0025_em-eta5-phi1*/	5,58,0,4,58,1,10,58,2,11,134,5,5,135,2,12,
/* out0026_em-eta6-phi1*/	5,57,0,3,57,1,13,58,2,4,134,4,6,134,5,11,
/* out0027_em-eta7-phi1*/	7,49,1,1,49,2,1,56,1,2,57,0,5,57,2,10,134,3,7,134,4,10,
/* out0028_em-eta8-phi1*/	5,49,2,2,56,0,8,56,1,6,56,2,1,134,3,9,
/* out0029_em-eta9-phi1*/	6,11,2,4,11,3,1,48,1,1,48,2,3,56,0,5,56,2,5,
/* out0030_em-eta10-phi1*/	5,11,2,12,11,3,3,11,4,9,11,5,12,48,2,1,
/* out0031_em-eta11-phi1*/	6,6,0,2,6,3,2,10,4,7,10,5,14,11,0,7,11,5,2,
/* out0032_em-eta12-phi1*/	4,6,0,13,6,1,1,9,2,9,10,4,5,
/* out0033_em-eta13-phi1*/	5,6,1,4,8,5,3,9,2,1,9,4,1,9,5,15,
/* out0034_em-eta14-phi1*/	4,2,0,1,2,3,6,8,4,2,8,5,10,
/* out0035_em-eta15-phi1*/	4,2,0,12,2,1,1,2,3,3,8,4,1,
/* out0036_em-eta16-phi1*/	4,2,0,2,2,1,9,5,2,1,5,5,2,
/* out0037_em-eta17-phi1*/	5,0,4,2,2,1,3,3,1,1,4,5,2,5,5,4,
/* out0038_em-eta18-phi1*/	4,0,4,6,0,5,8,1,0,1,4,5,1,
/* out0039_em-eta19-phi1*/	6,0,2,11,0,3,5,0,5,3,1,0,1,1,3,10,1,5,10,
/* out0040_em-eta0-phi2*/	1,141,0,16,
/* out0041_em-eta1-phi2*/	1,141,1,15,
/* out0042_em-eta2-phi2*/	4,70,1,4,140,0,16,140,1,1,141,1,1,
/* out0043_em-eta3-phi2*/	7,69,1,1,70,0,2,70,1,10,70,2,16,79,0,6,139,0,2,140,1,15,
/* out0044_em-eta4-phi2*/	6,69,0,8,69,1,14,69,2,9,79,0,1,139,0,14,139,1,4,
/* out0045_em-eta5-phi2*/	8,58,1,1,58,2,1,68,0,7,68,1,10,69,0,2,69,2,5,138,0,5,139,1,12,
/* out0046_em-eta6-phi2*/	7,57,1,3,57,2,1,67,1,2,68,0,9,68,2,6,138,0,11,138,1,6,
/* out0047_em-eta7-phi2*/	6,56,1,1,57,2,5,67,0,11,67,1,1,138,1,10,138,2,7,
/* out0048_em-eta8-phi2*/	5,56,1,7,56,2,4,66,0,1,67,0,3,138,2,9,
/* out0049_em-eta9-phi2*/	4,10,3,3,11,3,6,56,2,6,66,0,3,
/* out0050_em-eta10-phi2*/	6,10,0,1,10,1,1,10,2,11,10,3,13,11,3,6,11,4,7,
/* out0051_em-eta11-phi2*/	5,10,1,6,10,2,5,10,4,1,11,0,9,11,1,12,
/* out0052_em-eta12-phi2*/	5,9,2,6,9,3,14,9,4,2,10,4,3,11,1,3,
/* out0053_em-eta13-phi2*/	4,8,2,2,9,0,7,9,4,13,9,5,1,
/* out0054_em-eta14-phi2*/	4,8,4,6,8,5,3,9,0,7,9,1,3,
/* out0055_em-eta15-phi2*/	3,2,0,1,5,2,9,8,4,7,
/* out0056_em-eta16-phi2*/	3,5,2,5,5,4,2,5,5,6,
/* out0057_em-eta17-phi2*/	4,4,5,5,5,0,1,5,4,1,5,5,4,
/* out0058_em-eta18-phi2*/	3,0,5,2,4,4,3,4,5,6,
/* out0059_em-eta19-phi2*/	5,0,3,2,0,5,2,1,3,2,1,5,2,4,4,1,
/* out0060_em-eta0-phi3*/	1,141,3,16,
/* out0061_em-eta1-phi3*/	1,141,2,15,
/* out0062_em-eta2-phi3*/	3,140,2,1,140,3,16,141,2,1,
/* out0063_em-eta3-phi3*/	6,79,0,6,79,1,16,79,2,8,128,2,6,139,3,2,140,2,15,
/* out0064_em-eta4-phi3*/	8,69,1,1,69,2,2,78,0,7,78,1,10,79,0,3,79,2,7,139,2,4,139,3,14,
/* out0065_em-eta5-phi3*/	8,68,1,6,68,2,3,77,0,1,77,1,2,78,0,9,78,2,5,138,5,5,139,2,12,
/* out0066_em-eta6-phi3*/	5,67,1,5,68,2,7,77,0,9,138,4,6,138,5,11,
/* out0067_em-eta7-phi3*/	5,67,0,2,67,1,8,67,2,8,138,3,7,138,4,10,
/* out0068_em-eta8-phi3*/	4,66,0,1,66,1,7,67,2,6,138,3,9,
/* out0069_em-eta9-phi3*/	3,66,0,8,66,1,2,66,2,2,
/* out0070_em-eta10-phi3*/	4,10,0,13,13,2,9,66,0,3,66,2,2,
/* out0071_em-eta11-phi3*/	6,10,0,2,10,1,9,11,1,1,12,5,3,13,2,4,13,5,15,
/* out0072_em-eta12-phi3*/	6,8,0,3,8,2,1,8,3,14,9,3,2,12,4,1,12,5,8,
/* out0073_em-eta13-phi3*/	4,8,0,4,8,1,5,8,2,12,8,3,2,
/* out0074_em-eta14-phi3*/	4,8,1,6,8,2,1,9,0,2,9,1,11,
/* out0075_em-eta15-phi3*/	3,5,2,1,5,3,13,9,1,2,
/* out0076_em-eta16-phi3*/	3,4,2,1,5,3,2,5,4,11,
/* out0077_em-eta17-phi3*/	2,5,0,9,5,4,2,
/* out0078_em-eta18-phi3*/	4,4,4,5,4,5,2,5,0,2,5,1,1,
/* out0079_em-eta19-phi3*/	1,4,4,5,
/* out0080_em-eta0-phi4*/	1,145,0,16,
/* out0081_em-eta1-phi4*/	1,145,1,15,
/* out0082_em-eta2-phi4*/	6,128,1,5,128,2,5,129,0,3,144,0,16,144,1,1,145,1,1,
/* out0083_em-eta3-phi4*/	10,79,2,1,127,0,7,127,1,14,127,2,2,128,1,11,128,2,5,129,0,3,129,2,1,143,0,2,144,1,15,
/* out0084_em-eta4-phi4*/	8,78,1,6,78,2,4,126,0,3,126,1,3,127,0,9,127,2,7,143,0,14,143,1,4,
/* out0085_em-eta5-phi4*/	5,77,1,10,78,2,7,126,0,8,142,0,5,143,1,12,
/* out0086_em-eta6-phi4*/	5,77,0,5,77,1,4,77,2,12,142,0,11,142,1,6,
/* out0087_em-eta7-phi4*/	7,67,2,2,76,0,8,76,1,6,77,0,1,77,2,1,142,1,10,142,2,7,
/* out0088_em-eta8-phi4*/	3,66,1,6,76,0,8,142,2,9,
/* out0089_em-eta9-phi4*/	3,66,1,1,66,2,9,84,1,1,
/* out0090_em-eta10-phi4*/	6,12,2,1,12,3,6,13,2,3,13,3,16,13,4,2,66,2,3,
/* out0091_em-eta11-phi4*/	4,12,2,7,13,0,11,13,4,14,13,5,1,
/* out0092_em-eta12-phi4*/	5,8,0,1,12,4,14,12,5,5,13,0,4,13,1,3,
/* out0093_em-eta13-phi4*/	4,8,0,8,8,1,1,14,5,9,15,5,3,
/* out0094_em-eta14-phi4*/	3,8,1,4,14,4,11,14,5,2,
/* out0095_em-eta15-phi4*/	3,4,3,12,5,3,1,14,4,2,
/* out0096_em-eta16-phi4*/	2,4,2,9,4,3,4,
/* out0097_em-eta17-phi4*/	3,4,1,2,4,2,6,5,0,4,
/* out0098_em-eta18-phi4*/	1,5,1,9,
/* out0099_em-eta19-phi4*/	2,4,4,2,5,1,1,
/* out0100_em-eta0-phi5*/	1,145,3,16,
/* out0101_em-eta1-phi5*/	1,145,2,15,
/* out0102_em-eta2-phi5*/	4,129,0,3,144,2,1,144,3,16,145,2,1,
/* out0103_em-eta3-phi5*/	8,116,0,4,116,1,8,127,1,2,127,2,3,129,0,7,129,2,15,143,3,2,144,2,15,
/* out0104_em-eta4-phi5*/	6,116,0,12,126,1,12,126,2,2,127,2,4,143,2,4,143,3,14,
/* out0105_em-eta5-phi5*/	6,114,2,5,126,0,5,126,1,1,126,2,14,142,5,5,143,2,12,
/* out0106_em-eta6-phi5*/	6,76,1,1,77,2,3,114,1,14,114,2,3,142,4,6,142,5,11,
/* out0107_em-eta7-phi5*/	5,76,1,9,76,2,6,114,1,2,142,3,7,142,4,10,
/* out0108_em-eta8-phi5*/	3,76,2,10,84,2,5,142,3,9,
/* out0109_em-eta9-phi5*/	2,84,1,9,84,2,3,
/* out0110_em-eta10-phi5*/	3,12,0,7,12,3,9,84,1,6,
/* out0111_em-eta11-phi5*/	5,12,0,9,12,1,13,12,2,8,12,3,1,13,0,1,
/* out0112_em-eta12-phi5*/	5,12,1,3,12,4,1,13,1,13,15,2,7,15,5,3,
/* out0113_em-eta13-phi5*/	4,14,5,3,15,0,3,15,4,7,15,5,10,
/* out0114_em-eta14-phi5*/	4,14,4,2,14,5,2,15,0,12,15,1,3,
/* out0115_em-eta15-phi5*/	3,4,0,3,14,4,1,15,1,12,
/* out0116_em-eta16-phi5*/	2,4,0,12,4,1,1,
/* out0117_em-eta17-phi5*/	2,4,0,1,4,1,10,
/* out0118_em-eta18-phi5*/	2,4,1,3,5,1,5,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	1,149,0,16,
/* out0121_em-eta1-phi6*/	1,149,1,15,
/* out0122_em-eta2-phi6*/	4,118,2,3,148,0,16,148,1,1,149,1,1,
/* out0123_em-eta3-phi6*/	8,116,1,8,116,2,4,117,1,3,117,2,2,118,0,15,118,2,7,147,0,2,148,1,15,
/* out0124_em-eta4-phi6*/	6,115,1,2,115,2,12,116,2,12,117,1,4,147,0,14,147,1,4,
/* out0125_em-eta5-phi6*/	6,114,2,5,115,0,5,115,1,14,115,2,1,146,0,5,147,1,12,
/* out0126_em-eta6-phi6*/	6,85,2,1,86,1,3,114,0,14,114,2,3,146,0,11,146,1,6,
/* out0127_em-eta7-phi6*/	5,85,1,7,85,2,9,114,0,2,146,1,10,146,2,7,
/* out0128_em-eta8-phi6*/	3,84,2,5,85,1,9,146,2,9,
/* out0129_em-eta9-phi6*/	2,84,0,9,84,2,3,
/* out0130_em-eta10-phi6*/	4,16,5,1,17,2,3,17,5,12,84,0,6,
/* out0131_em-eta11-phi6*/	5,16,4,5,16,5,15,17,0,7,17,4,2,17,5,2,
/* out0132_em-eta12-phi6*/	4,15,2,8,15,3,3,16,4,11,17,1,6,
/* out0133_em-eta13-phi6*/	5,14,2,3,14,3,2,15,2,1,15,3,9,15,4,9,
/* out0134_em-eta14-phi6*/	5,14,0,1,14,1,4,14,2,13,14,3,1,15,0,1,
/* out0135_em-eta15-phi6*/	3,14,1,12,15,1,1,19,5,3,
/* out0136_em-eta16-phi6*/	2,18,5,8,19,5,5,
/* out0137_em-eta17-phi6*/	2,18,4,5,18,5,6,
/* out0138_em-eta18-phi6*/	1,18,4,8,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	1,149,3,16,
/* out0141_em-eta1-phi7*/	1,149,2,15,
/* out0142_em-eta2-phi7*/	6,118,2,3,119,0,5,119,1,5,148,2,1,148,3,16,149,2,1,
/* out0143_em-eta3-phi7*/	10,88,1,1,117,0,7,117,1,2,117,2,14,118,0,1,118,2,3,119,0,5,119,1,11,147,3,2,148,2,15,
/* out0144_em-eta4-phi7*/	8,87,1,4,87,2,6,115,0,3,115,2,3,117,0,9,117,1,7,147,2,4,147,3,14,
/* out0145_em-eta5-phi7*/	5,86,2,10,87,1,7,115,0,8,146,5,5,147,2,12,
/* out0146_em-eta6-phi7*/	5,86,0,5,86,1,12,86,2,4,146,4,6,146,5,11,
/* out0147_em-eta7-phi7*/	7,85,0,8,85,2,6,86,0,1,86,1,1,95,1,2,146,3,7,146,4,10,
/* out0148_em-eta8-phi7*/	3,85,0,8,94,2,6,146,3,9,
/* out0149_em-eta9-phi7*/	3,84,0,1,94,1,9,94,2,1,
/* out0150_em-eta10-phi7*/	5,17,2,13,17,3,11,17,4,3,17,5,2,94,1,3,
/* out0151_em-eta11-phi7*/	5,16,1,1,16,2,14,16,3,1,17,0,7,17,4,11,
/* out0152_em-eta12-phi7*/	6,15,3,1,16,1,12,16,2,2,17,0,2,17,1,10,21,5,1,
/* out0153_em-eta13-phi7*/	4,14,3,10,15,3,3,20,5,7,21,5,2,
/* out0154_em-eta14-phi7*/	3,14,0,12,14,3,3,20,4,5,
/* out0155_em-eta15-phi7*/	3,14,0,3,19,2,10,19,5,4,
/* out0156_em-eta16-phi7*/	3,19,0,2,19,4,7,19,5,4,
/* out0157_em-eta17-phi7*/	2,18,5,2,19,0,9,
/* out0158_em-eta18-phi7*/	3,18,4,3,19,0,1,19,1,6,
/* out0159_em-eta19-phi7*/	1,19,1,2,
/* out0160_em-eta0-phi8*/	1,153,0,16,
/* out0161_em-eta1-phi8*/	1,153,1,15,
/* out0162_em-eta2-phi8*/	3,152,0,16,152,1,1,153,1,1,
/* out0163_em-eta3-phi8*/	6,88,0,6,88,1,8,88,2,16,119,0,6,151,0,2,152,1,15,
/* out0164_em-eta4-phi8*/	8,87,0,7,87,2,10,88,0,3,88,1,7,97,1,2,97,2,1,151,0,14,151,1,4,
/* out0165_em-eta5-phi8*/	8,86,0,1,86,2,2,87,0,9,87,1,5,96,1,3,96,2,6,150,0,5,151,1,12,
/* out0166_em-eta6-phi8*/	5,86,0,9,95,2,5,96,1,7,150,0,11,150,1,6,
/* out0167_em-eta7-phi8*/	5,95,0,2,95,1,8,95,2,8,150,1,10,150,2,7,
/* out0168_em-eta8-phi8*/	4,94,0,1,94,2,7,95,1,6,150,2,9,
/* out0169_em-eta9-phi8*/	3,94,0,8,94,1,2,94,2,2,
/* out0170_em-eta10-phi8*/	6,16,3,4,17,3,5,22,5,6,23,5,7,94,0,3,94,1,2,
/* out0171_em-eta11-phi8*/	4,16,0,10,16,3,11,22,4,7,22,5,5,
/* out0172_em-eta12-phi8*/	5,16,0,6,16,1,3,21,2,10,21,4,1,21,5,8,
/* out0173_em-eta13-phi8*/	4,20,5,7,21,0,7,21,4,5,21,5,5,
/* out0174_em-eta14-phi8*/	4,20,4,10,20,5,2,21,0,3,21,1,4,
/* out0175_em-eta15-phi8*/	4,19,2,6,19,3,7,20,4,1,21,1,1,
/* out0176_em-eta16-phi8*/	3,18,2,3,19,3,2,19,4,9,
/* out0177_em-eta17-phi8*/	2,18,2,8,19,0,3,
/* out0178_em-eta18-phi8*/	4,18,1,4,18,2,1,19,0,1,19,1,4,
/* out0179_em-eta19-phi8*/	2,18,1,2,19,1,4,
/* out0180_em-eta0-phi9*/	1,153,3,16,
/* out0181_em-eta1-phi9*/	1,153,2,15,
/* out0182_em-eta2-phi9*/	4,98,2,4,152,2,1,152,3,16,153,2,1,
/* out0183_em-eta3-phi9*/	7,88,0,6,97,2,1,98,0,2,98,1,16,98,2,10,151,3,2,152,2,15,
/* out0184_em-eta4-phi9*/	6,88,0,1,97,0,8,97,1,9,97,2,14,151,2,4,151,3,14,
/* out0185_em-eta5-phi9*/	8,96,0,7,96,2,10,97,0,2,97,1,5,106,1,1,106,2,1,150,5,5,151,2,12,
/* out0186_em-eta6-phi9*/	7,95,2,2,96,0,9,96,1,6,105,1,1,105,2,3,150,4,6,150,5,11,
/* out0187_em-eta7-phi9*/	6,95,0,11,95,2,1,104,2,1,105,1,5,150,3,7,150,4,10,
/* out0188_em-eta8-phi9*/	5,94,0,1,95,0,3,104,1,4,104,2,7,150,3,9,
/* out0189_em-eta9-phi9*/	3,23,2,8,94,0,3,104,1,6,
/* out0190_em-eta10-phi9*/	7,22,2,1,22,5,1,23,0,3,23,2,8,23,3,4,23,4,14,23,5,9,
/* out0191_em-eta11-phi9*/	5,22,2,1,22,4,7,22,5,4,23,0,13,23,1,8,
/* out0192_em-eta12-phi9*/	6,20,3,1,21,2,6,21,3,14,21,4,2,22,4,2,23,1,3,
/* out0193_em-eta13-phi9*/	4,20,2,12,20,3,1,21,0,2,21,4,8,
/* out0194_em-eta14-phi9*/	4,20,1,7,20,2,3,21,0,4,21,1,6,
/* out0195_em-eta15-phi9*/	4,18,3,3,19,3,6,20,1,2,21,1,5,
/* out0196_em-eta16-phi9*/	3,18,2,1,18,3,11,19,3,1,
/* out0197_em-eta17-phi9*/	4,18,0,5,18,1,2,18,2,3,18,3,1,
/* out0198_em-eta18-phi9*/	3,18,0,2,18,1,7,24,3,1,
/* out0199_em-eta19-phi9*/	5,18,1,1,24,3,2,24,5,1,25,3,2,25,5,2,
/* out0200_em-eta0-phi10*/	1,157,0,16,
/* out0201_em-eta1-phi10*/	1,157,1,15,
/* out0202_em-eta2-phi10*/	6,98,2,1,108,0,1,108,1,1,156,0,16,156,1,1,157,1,1,
/* out0203_em-eta3-phi10*/	7,98,0,14,98,2,1,107,2,11,108,0,3,108,1,13,155,0,2,156,1,15,
/* out0204_em-eta4-phi10*/	7,97,0,6,106,2,5,107,0,2,107,1,15,107,2,3,155,0,14,155,1,4,
/* out0205_em-eta5-phi10*/	5,106,0,4,106,1,11,106,2,10,154,0,5,155,1,12,
/* out0206_em-eta6-phi10*/	5,105,0,3,105,2,13,106,1,4,154,0,11,154,1,6,
/* out0207_em-eta7-phi10*/	5,104,2,2,105,0,5,105,1,10,154,1,10,154,2,7,
/* out0208_em-eta8-phi10*/	4,104,0,8,104,1,1,104,2,6,154,2,9,
/* out0209_em-eta9-phi10*/	4,23,3,4,52,0,1,104,0,5,104,1,5,
/* out0210_em-eta10-phi10*/	6,22,0,4,22,2,7,22,3,16,23,3,8,23,4,2,52,0,1,
/* out0211_em-eta11-phi10*/	5,22,0,8,22,1,14,22,2,7,23,1,2,31,5,2,
/* out0212_em-eta12-phi10*/	6,20,3,6,21,3,2,22,1,2,23,1,3,30,5,8,31,5,5,
/* out0213_em-eta13-phi10*/	5,20,0,11,20,2,1,20,3,8,30,4,2,30,5,1,
/* out0214_em-eta14-phi10*/	4,20,0,5,20,1,7,29,2,3,29,5,3,
/* out0215_em-eta15-phi10*/	2,28,5,7,29,5,9,
/* out0216_em-eta16-phi10*/	4,18,0,2,18,3,1,28,4,3,28,5,7,
/* out0217_em-eta17-phi10*/	3,18,0,6,24,0,2,28,4,3,
/* out0218_em-eta18-phi10*/	3,18,0,1,24,0,5,24,3,8,
/* out0219_em-eta19-phi10*/	5,24,2,1,24,3,3,24,5,5,25,3,9,25,5,9,
/* out0220_em-eta0-phi11*/	1,157,3,16,
/* out0221_em-eta1-phi11*/	1,157,2,15,
/* out0222_em-eta2-phi11*/	3,156,2,1,156,3,16,157,2,1,
/* out0223_em-eta3-phi11*/	6,107,0,4,107,2,2,108,0,12,108,1,2,155,3,2,156,2,15,
/* out0224_em-eta4-phi11*/	7,55,0,11,55,1,4,106,0,1,107,0,10,107,1,1,155,2,4,155,3,14,
/* out0225_em-eta5-phi11*/	7,54,0,3,54,1,3,55,0,5,55,2,4,106,0,10,154,5,5,155,2,12,
/* out0226_em-eta6-phi11*/	7,54,0,13,54,1,1,54,2,3,105,0,4,106,0,1,154,4,6,154,5,11,
/* out0227_em-eta7-phi11*/	6,53,0,9,53,1,4,54,2,1,105,0,4,154,3,7,154,4,10,
/* out0228_em-eta8-phi11*/	4,53,0,7,53,2,4,104,0,2,154,3,9,
/* out0229_em-eta9-phi11*/	3,52,0,8,52,1,3,104,0,1,
/* out0230_em-eta10-phi11*/	3,22,0,1,52,0,6,52,2,3,
/* out0231_em-eta11-phi11*/	6,22,0,3,31,2,16,31,3,4,31,4,3,31,5,4,52,2,1,
/* out0232_em-eta12-phi11*/	4,30,5,5,31,0,9,31,4,9,31,5,5,
/* out0233_em-eta13-phi11*/	5,29,2,1,30,4,14,30,5,2,31,0,2,31,1,4,
/* out0234_em-eta14-phi11*/	4,29,2,12,29,3,4,29,4,2,29,5,2,
/* out0235_em-eta15-phi11*/	3,29,0,5,29,4,9,29,5,2,
/* out0236_em-eta16-phi11*/	4,28,4,3,28,5,2,29,0,6,29,1,2,
/* out0237_em-eta17-phi11*/	3,24,0,5,28,4,7,29,1,2,
/* out0238_em-eta18-phi11*/	4,24,0,4,24,1,3,24,2,9,24,3,2,
/* out0239_em-eta19-phi11*/	5,24,2,1,24,5,8,25,0,4,25,3,5,25,5,5,
/* out0240_em-eta0-phi12*/	1,161,0,16,
/* out0241_em-eta1-phi12*/	1,161,1,15,
/* out0242_em-eta2-phi12*/	3,160,0,16,160,1,1,161,1,1,
/* out0243_em-eta3-phi12*/	6,64,0,4,64,1,2,65,0,12,65,2,2,159,0,2,160,1,15,
/* out0244_em-eta4-phi12*/	7,55,1,12,55,2,4,63,0,1,64,0,10,64,2,1,159,0,14,159,1,4,
/* out0245_em-eta5-phi12*/	5,54,1,7,55,2,8,63,0,10,158,0,5,159,1,12,
/* out0246_em-eta6-phi12*/	6,54,1,5,54,2,11,62,0,4,63,0,1,158,0,11,158,1,6,
/* out0247_em-eta7-phi12*/	6,53,1,12,53,2,1,54,2,1,62,0,4,158,1,10,158,2,7,
/* out0248_em-eta8-phi12*/	4,52,1,1,53,2,11,61,0,2,158,2,9,
/* out0249_em-eta9-phi12*/	2,52,1,11,61,0,1,
/* out0250_em-eta10-phi12*/	2,37,5,1,52,2,10,
/* out0251_em-eta11-phi12*/	7,30,2,1,30,3,11,31,3,12,31,4,2,36,5,2,37,5,1,52,2,1,
/* out0252_em-eta12-phi12*/	6,30,0,1,30,1,4,30,2,15,30,3,3,31,0,3,31,4,2,
/* out0253_em-eta13-phi12*/	4,29,3,1,30,1,7,31,0,2,31,1,12,
/* out0254_em-eta14-phi12*/	4,28,2,1,28,3,6,29,3,11,29,4,2,
/* out0255_em-eta15-phi12*/	4,28,2,12,28,3,1,29,0,1,29,4,3,
/* out0256_em-eta16-phi12*/	4,28,1,3,28,2,3,29,0,4,29,1,3,
/* out0257_em-eta17-phi12*/	2,24,1,6,29,1,8,
/* out0258_em-eta18-phi12*/	5,24,1,6,24,2,5,24,4,1,25,0,12,25,1,5,
/* out0259_em-eta19-phi12*/	2,24,4,4,24,5,2,
/* out0260_em-eta0-phi13*/	1,161,3,16,
/* out0261_em-eta1-phi13*/	1,161,2,15,
/* out0262_em-eta2-phi13*/	6,65,0,1,65,2,1,75,1,1,160,2,1,160,3,16,161,2,1,
/* out0263_em-eta3-phi13*/	7,64,1,11,65,0,3,65,2,13,75,0,14,75,1,1,159,3,2,160,2,15,
/* out0264_em-eta4-phi13*/	7,63,1,5,64,0,2,64,1,3,64,2,15,74,0,6,159,2,4,159,3,14,
/* out0265_em-eta5-phi13*/	5,63,0,4,63,1,10,63,2,11,158,5,5,159,2,12,
/* out0266_em-eta6-phi13*/	5,62,0,3,62,1,13,63,2,4,158,4,6,158,5,11,
/* out0267_em-eta7-phi13*/	5,61,1,2,62,0,5,62,2,10,158,3,7,158,4,10,
/* out0268_em-eta8-phi13*/	4,61,0,8,61,1,6,61,2,1,158,3,9,
/* out0269_em-eta9-phi13*/	5,37,2,4,37,3,1,52,1,1,61,0,5,61,2,5,
/* out0270_em-eta10-phi13*/	5,37,2,12,37,3,3,37,4,9,37,5,12,52,2,1,
/* out0271_em-eta11-phi13*/	6,30,0,2,30,3,2,36,4,7,36,5,14,37,0,7,37,5,2,
/* out0272_em-eta12-phi13*/	4,30,0,13,30,1,1,33,2,9,36,4,5,
/* out0273_em-eta13-phi13*/	5,30,1,4,32,5,3,33,2,1,33,4,1,33,5,15,
/* out0274_em-eta14-phi13*/	4,28,0,1,28,3,6,32,4,2,32,5,10,
/* out0275_em-eta15-phi13*/	4,28,0,12,28,1,1,28,3,3,32,4,1,
/* out0276_em-eta16-phi13*/	4,27,2,1,27,5,2,28,0,2,28,1,9,
/* out0277_em-eta17-phi13*/	6,24,1,1,25,1,2,26,5,2,27,5,4,28,1,3,29,1,1,
/* out0278_em-eta18-phi13*/	3,24,4,3,25,1,9,26,5,1,
/* out0279_em-eta19-phi13*/	1,24,4,5,
/* out0280_em-eta0-phi14*/	1,165,0,16,
/* out0281_em-eta1-phi14*/	1,165,1,15,
/* out0282_em-eta2-phi14*/	4,75,1,4,164,0,16,164,1,1,165,1,1,
/* out0283_em-eta3-phi14*/	7,74,1,1,75,0,2,75,1,10,75,2,16,83,0,6,163,0,2,164,1,15,
/* out0284_em-eta4-phi14*/	6,74,0,8,74,1,14,74,2,9,83,0,1,163,0,14,163,1,4,
/* out0285_em-eta5-phi14*/	8,63,1,1,63,2,1,73,0,7,73,1,10,74,0,2,74,2,5,162,0,5,163,1,12,
/* out0286_em-eta6-phi14*/	7,62,1,3,62,2,1,72,1,2,73,0,9,73,2,6,162,0,11,162,1,6,
/* out0287_em-eta7-phi14*/	6,61,1,1,62,2,5,72,0,11,72,1,1,162,1,10,162,2,7,
/* out0288_em-eta8-phi14*/	5,61,1,7,61,2,4,71,0,1,72,0,3,162,2,9,
/* out0289_em-eta9-phi14*/	4,36,3,3,37,3,6,61,2,6,71,0,3,
/* out0290_em-eta10-phi14*/	6,36,0,1,36,1,1,36,2,11,36,3,13,37,3,6,37,4,7,
/* out0291_em-eta11-phi14*/	5,36,1,6,36,2,5,36,4,1,37,0,9,37,1,12,
/* out0292_em-eta12-phi14*/	5,33,2,6,33,3,14,33,4,2,36,4,3,37,1,3,
/* out0293_em-eta13-phi14*/	4,32,2,2,33,0,7,33,4,13,33,5,1,
/* out0294_em-eta14-phi14*/	4,32,4,6,32,5,3,33,0,7,33,1,3,
/* out0295_em-eta15-phi14*/	3,27,2,9,28,0,1,32,4,7,
/* out0296_em-eta16-phi14*/	3,27,2,5,27,4,2,27,5,6,
/* out0297_em-eta17-phi14*/	4,26,5,5,27,0,1,27,4,1,27,5,4,
/* out0298_em-eta18-phi14*/	3,24,4,1,26,4,3,26,5,6,
/* out0299_em-eta19-phi14*/	2,24,4,2,26,4,1,
/* out0300_em-eta0-phi15*/	1,165,3,16,
/* out0301_em-eta1-phi15*/	1,165,2,15,
/* out0302_em-eta2-phi15*/	3,164,2,1,164,3,16,165,2,1,
/* out0303_em-eta3-phi15*/	6,83,0,6,83,1,16,83,2,8,133,0,6,163,3,2,164,2,15,
/* out0304_em-eta4-phi15*/	8,74,1,1,74,2,2,82,0,7,82,1,10,83,0,3,83,2,7,163,2,4,163,3,14,
/* out0305_em-eta5-phi15*/	8,73,1,6,73,2,3,81,0,1,81,1,2,82,0,9,82,2,5,162,5,5,163,2,12,
/* out0306_em-eta6-phi15*/	5,72,1,5,73,2,7,81,0,9,162,4,6,162,5,11,
/* out0307_em-eta7-phi15*/	5,72,0,2,72,1,8,72,2,8,162,3,7,162,4,10,
/* out0308_em-eta8-phi15*/	4,71,0,1,71,1,7,72,2,6,162,3,9,
/* out0309_em-eta9-phi15*/	3,71,0,8,71,1,2,71,2,2,
/* out0310_em-eta10-phi15*/	4,35,2,9,36,0,13,71,0,3,71,2,2,
/* out0311_em-eta11-phi15*/	6,34,5,3,35,2,4,35,5,15,36,0,2,36,1,9,37,1,1,
/* out0312_em-eta12-phi15*/	6,32,0,3,32,2,1,32,3,14,33,3,2,34,4,1,34,5,8,
/* out0313_em-eta13-phi15*/	4,32,0,4,32,1,5,32,2,12,32,3,2,
/* out0314_em-eta14-phi15*/	4,32,1,6,32,2,1,33,0,2,33,1,11,
/* out0315_em-eta15-phi15*/	3,27,2,1,27,3,13,33,1,2,
/* out0316_em-eta16-phi15*/	3,26,2,1,27,3,2,27,4,11,
/* out0317_em-eta17-phi15*/	2,27,0,9,27,4,2,
/* out0318_em-eta18-phi15*/	4,26,4,5,26,5,2,27,0,2,27,1,1,
/* out0319_em-eta19-phi15*/	1,26,4,5,
/* out0320_em-eta0-phi16*/	1,169,0,16,
/* out0321_em-eta1-phi16*/	1,169,1,15,
/* out0322_em-eta2-phi16*/	6,132,0,3,133,0,5,133,2,5,168,0,16,168,1,1,169,1,1,
/* out0323_em-eta3-phi16*/	10,83,2,1,131,0,7,131,1,14,131,2,2,132,0,3,132,2,1,133,0,5,133,2,11,167,0,2,168,1,15,
/* out0324_em-eta4-phi16*/	8,82,1,6,82,2,4,130,0,3,130,1,3,131,0,9,131,2,7,167,0,14,167,1,4,
/* out0325_em-eta5-phi16*/	5,81,1,10,82,2,7,130,0,8,166,0,5,167,1,12,
/* out0326_em-eta6-phi16*/	5,81,0,5,81,1,4,81,2,12,166,0,11,166,1,6,
/* out0327_em-eta7-phi16*/	7,72,2,2,80,0,8,80,1,6,81,0,1,81,2,1,166,1,10,166,2,7,
/* out0328_em-eta8-phi16*/	3,71,1,6,80,0,8,166,2,9,
/* out0329_em-eta9-phi16*/	3,71,1,1,71,2,9,89,1,1,
/* out0330_em-eta10-phi16*/	6,34,2,1,34,3,6,35,2,3,35,3,16,35,4,2,71,2,3,
/* out0331_em-eta11-phi16*/	4,34,2,7,35,0,11,35,4,14,35,5,1,
/* out0332_em-eta12-phi16*/	5,32,0,1,34,4,14,34,5,5,35,0,4,35,1,3,
/* out0333_em-eta13-phi16*/	4,32,0,8,32,1,1,38,5,9,39,5,3,
/* out0334_em-eta14-phi16*/	3,32,1,4,38,4,11,38,5,2,
/* out0335_em-eta15-phi16*/	3,26,3,12,27,3,1,38,4,2,
/* out0336_em-eta16-phi16*/	2,26,2,9,26,3,4,
/* out0337_em-eta17-phi16*/	3,26,1,2,26,2,6,27,0,4,
/* out0338_em-eta18-phi16*/	1,27,1,9,
/* out0339_em-eta19-phi16*/	2,26,4,2,27,1,1,
/* out0340_em-eta0-phi17*/	1,169,3,16,
/* out0341_em-eta1-phi17*/	1,169,2,15,
/* out0342_em-eta2-phi17*/	4,132,0,3,168,2,1,168,3,16,169,2,1,
/* out0343_em-eta3-phi17*/	8,124,0,4,124,1,8,131,1,2,131,2,3,132,0,7,132,2,15,167,3,2,168,2,15,
/* out0344_em-eta4-phi17*/	6,124,0,12,130,1,12,130,2,2,131,2,4,167,2,4,167,3,14,
/* out0345_em-eta5-phi17*/	6,120,2,5,130,0,5,130,1,1,130,2,14,166,5,5,167,2,12,
/* out0346_em-eta6-phi17*/	6,80,1,1,81,2,3,120,1,14,120,2,3,166,4,6,166,5,11,
/* out0347_em-eta7-phi17*/	5,80,1,9,80,2,7,120,1,2,166,3,7,166,4,10,
/* out0348_em-eta8-phi17*/	3,80,2,9,89,2,4,166,3,9,
/* out0349_em-eta9-phi17*/	2,89,1,9,89,2,3,
/* out0350_em-eta10-phi17*/	3,34,0,7,34,3,9,89,1,6,
/* out0351_em-eta11-phi17*/	5,34,0,9,34,1,13,34,2,8,34,3,1,35,0,1,
/* out0352_em-eta12-phi17*/	5,34,1,3,34,4,1,35,1,13,39,2,7,39,5,3,
/* out0353_em-eta13-phi17*/	4,38,5,3,39,0,3,39,4,7,39,5,10,
/* out0354_em-eta14-phi17*/	4,38,4,2,38,5,2,39,0,12,39,1,3,
/* out0355_em-eta15-phi17*/	3,26,0,3,38,4,1,39,1,12,
/* out0356_em-eta16-phi17*/	2,26,0,12,26,1,1,
/* out0357_em-eta17-phi17*/	2,26,0,1,26,1,10,
/* out0358_em-eta18-phi17*/	2,26,1,3,27,1,5,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	1,173,0,16,
/* out0361_em-eta1-phi18*/	1,173,1,15,
/* out0362_em-eta2-phi18*/	4,125,0,3,172,0,16,172,1,1,173,1,1,
/* out0363_em-eta3-phi18*/	8,122,1,3,122,2,2,124,1,8,124,2,4,125,0,7,125,1,15,171,0,2,172,1,15,
/* out0364_em-eta4-phi18*/	6,121,1,2,121,2,12,122,1,4,124,2,12,171,0,14,171,1,4,
/* out0365_em-eta5-phi18*/	6,120,2,5,121,0,5,121,1,14,121,2,1,170,0,5,171,1,12,
/* out0366_em-eta6-phi18*/	6,90,2,1,91,1,3,120,0,14,120,2,3,170,0,11,170,1,6,
/* out0367_em-eta7-phi18*/	5,90,1,7,90,2,9,120,0,2,170,1,10,170,2,7,
/* out0368_em-eta8-phi18*/	3,89,2,5,90,1,9,170,2,9,
/* out0369_em-eta9-phi18*/	2,89,0,9,89,2,4,
/* out0370_em-eta10-phi18*/	4,40,5,1,41,2,3,41,5,12,89,0,6,
/* out0371_em-eta11-phi18*/	5,40,4,5,40,5,15,41,0,7,41,4,2,41,5,2,
/* out0372_em-eta12-phi18*/	4,39,2,8,39,3,3,40,4,11,41,1,6,
/* out0373_em-eta13-phi18*/	5,38,2,3,38,3,2,39,2,1,39,3,9,39,4,9,
/* out0374_em-eta14-phi18*/	5,38,0,1,38,1,4,38,2,13,38,3,1,39,0,1,
/* out0375_em-eta15-phi18*/	3,38,1,12,39,1,1,43,5,3,
/* out0376_em-eta16-phi18*/	2,42,5,8,43,5,5,
/* out0377_em-eta17-phi18*/	2,42,4,5,42,5,6,
/* out0378_em-eta18-phi18*/	1,42,4,8,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	1,173,3,16,
/* out0381_em-eta1-phi19*/	1,173,2,15,
/* out0382_em-eta2-phi19*/	6,123,0,5,123,1,5,125,0,3,172,2,1,172,3,16,173,2,1,
/* out0383_em-eta3-phi19*/	10,93,1,1,122,0,7,122,1,2,122,2,14,123,0,5,123,1,11,125,0,3,125,1,1,171,3,2,172,2,15,
/* out0384_em-eta4-phi19*/	8,92,1,4,92,2,6,121,0,3,121,2,3,122,0,9,122,1,7,171,2,4,171,3,14,
/* out0385_em-eta5-phi19*/	5,91,2,10,92,1,7,121,0,8,170,5,5,171,2,12,
/* out0386_em-eta6-phi19*/	5,91,0,5,91,1,12,91,2,4,170,4,6,170,5,11,
/* out0387_em-eta7-phi19*/	7,90,0,8,90,2,6,91,0,1,91,1,1,100,1,2,170,3,7,170,4,10,
/* out0388_em-eta8-phi19*/	3,90,0,8,99,2,6,170,3,9,
/* out0389_em-eta9-phi19*/	3,89,0,1,99,1,9,99,2,1,
/* out0390_em-eta10-phi19*/	5,41,2,13,41,3,11,41,4,3,41,5,2,99,1,3,
/* out0391_em-eta11-phi19*/	5,40,1,1,40,2,14,40,3,1,41,0,7,41,4,11,
/* out0392_em-eta12-phi19*/	6,39,3,1,40,1,12,40,2,2,41,0,2,41,1,10,45,5,1,
/* out0393_em-eta13-phi19*/	4,38,3,10,39,3,3,44,5,7,45,5,2,
/* out0394_em-eta14-phi19*/	3,38,0,12,38,3,3,44,4,5,
/* out0395_em-eta15-phi19*/	3,38,0,3,43,2,10,43,5,4,
/* out0396_em-eta16-phi19*/	3,43,0,2,43,4,7,43,5,4,
/* out0397_em-eta17-phi19*/	2,42,5,2,43,0,9,
/* out0398_em-eta18-phi19*/	3,42,4,3,43,0,1,43,1,6,
/* out0399_em-eta19-phi19*/	1,43,1,2,
/* out0400_em-eta0-phi20*/	1,177,0,16,
/* out0401_em-eta1-phi20*/	1,177,1,15,
/* out0402_em-eta2-phi20*/	3,176,0,16,176,1,1,177,1,1,
/* out0403_em-eta3-phi20*/	6,93,0,6,93,1,8,93,2,16,123,0,6,175,0,2,176,1,15,
/* out0404_em-eta4-phi20*/	8,92,0,7,92,2,10,93,0,3,93,1,7,102,1,2,102,2,1,175,0,14,175,1,4,
/* out0405_em-eta5-phi20*/	8,91,0,1,91,2,2,92,0,9,92,1,5,101,1,3,101,2,6,174,0,5,175,1,12,
/* out0406_em-eta6-phi20*/	5,91,0,9,100,2,5,101,1,7,174,0,11,174,1,6,
/* out0407_em-eta7-phi20*/	5,100,0,2,100,1,8,100,2,8,174,1,10,174,2,7,
/* out0408_em-eta8-phi20*/	4,99,0,1,99,2,7,100,1,6,174,2,9,
/* out0409_em-eta9-phi20*/	3,99,0,8,99,1,2,99,2,2,
/* out0410_em-eta10-phi20*/	6,40,3,4,41,3,5,46,5,6,47,5,7,99,0,3,99,1,2,
/* out0411_em-eta11-phi20*/	4,40,0,10,40,3,11,46,4,7,46,5,5,
/* out0412_em-eta12-phi20*/	5,40,0,6,40,1,3,45,2,10,45,4,1,45,5,8,
/* out0413_em-eta13-phi20*/	4,44,5,7,45,0,7,45,4,5,45,5,5,
/* out0414_em-eta14-phi20*/	4,44,4,10,44,5,2,45,0,3,45,1,4,
/* out0415_em-eta15-phi20*/	4,43,2,6,43,3,7,44,4,1,45,1,1,
/* out0416_em-eta16-phi20*/	3,42,2,3,43,3,2,43,4,9,
/* out0417_em-eta17-phi20*/	2,42,2,8,43,0,3,
/* out0418_em-eta18-phi20*/	4,42,1,4,42,2,1,43,0,1,43,1,4,
/* out0419_em-eta19-phi20*/	2,42,1,2,43,1,4,
/* out0420_em-eta0-phi21*/	1,177,3,16,
/* out0421_em-eta1-phi21*/	1,177,2,15,
/* out0422_em-eta2-phi21*/	4,103,2,4,176,2,1,176,3,16,177,2,1,
/* out0423_em-eta3-phi21*/	7,93,0,6,102,2,1,103,0,2,103,1,16,103,2,10,175,3,2,176,2,15,
/* out0424_em-eta4-phi21*/	6,93,0,1,102,0,8,102,1,9,102,2,14,175,2,4,175,3,14,
/* out0425_em-eta5-phi21*/	8,101,0,7,101,2,10,102,0,2,102,1,5,111,1,1,111,2,1,174,5,5,175,2,12,
/* out0426_em-eta6-phi21*/	7,100,2,2,101,0,9,101,1,6,110,1,1,110,2,3,174,4,6,174,5,11,
/* out0427_em-eta7-phi21*/	6,100,0,11,100,2,1,109,2,1,110,1,5,174,3,7,174,4,10,
/* out0428_em-eta8-phi21*/	5,99,0,1,100,0,3,109,1,4,109,2,7,174,3,9,
/* out0429_em-eta9-phi21*/	3,47,2,8,99,0,3,109,1,6,
/* out0430_em-eta10-phi21*/	7,46,2,1,46,5,1,47,0,3,47,2,8,47,3,4,47,4,14,47,5,9,
/* out0431_em-eta11-phi21*/	5,46,2,1,46,4,7,46,5,4,47,0,13,47,1,8,
/* out0432_em-eta12-phi21*/	6,44,3,1,45,2,6,45,3,14,45,4,2,46,4,2,47,1,3,
/* out0433_em-eta13-phi21*/	4,44,2,12,44,3,1,45,0,2,45,4,8,
/* out0434_em-eta14-phi21*/	4,44,1,7,44,2,3,45,0,4,45,1,6,
/* out0435_em-eta15-phi21*/	4,42,3,3,43,3,6,44,1,2,45,1,5,
/* out0436_em-eta16-phi21*/	3,42,2,1,42,3,11,43,3,1,
/* out0437_em-eta17-phi21*/	4,42,0,5,42,1,2,42,2,3,42,3,1,
/* out0438_em-eta18-phi21*/	2,42,0,2,42,1,7,
/* out0439_em-eta19-phi21*/	1,42,1,1,
/* out0440_em-eta0-phi22*/	1,181,0,16,
/* out0441_em-eta1-phi22*/	1,181,1,15,
/* out0442_em-eta2-phi22*/	6,103,2,1,113,0,1,113,1,1,180,0,16,180,1,1,181,1,1,
/* out0443_em-eta3-phi22*/	7,103,0,14,103,2,1,112,2,11,113,0,3,113,1,13,179,0,2,180,1,15,
/* out0444_em-eta4-phi22*/	7,102,0,6,111,2,5,112,0,2,112,1,15,112,2,3,179,0,14,179,1,4,
/* out0445_em-eta5-phi22*/	5,111,0,4,111,1,11,111,2,10,178,0,5,179,1,12,
/* out0446_em-eta6-phi22*/	5,110,0,3,110,2,13,111,1,4,178,0,11,178,1,6,
/* out0447_em-eta7-phi22*/	5,109,2,2,110,0,5,110,1,10,178,1,10,178,2,7,
/* out0448_em-eta8-phi22*/	4,109,0,8,109,1,1,109,2,6,178,2,9,
/* out0449_em-eta9-phi22*/	3,47,3,4,109,0,5,109,1,5,
/* out0450_em-eta10-phi22*/	5,46,0,4,46,2,7,46,3,16,47,3,8,47,4,2,
/* out0451_em-eta11-phi22*/	4,46,0,8,46,1,14,46,2,7,47,1,2,
/* out0452_em-eta12-phi22*/	4,44,3,6,45,3,2,46,1,2,47,1,3,
/* out0453_em-eta13-phi22*/	3,44,0,11,44,2,1,44,3,8,
/* out0454_em-eta14-phi22*/	2,44,0,5,44,1,7,
/* out0455_em-eta15-phi22*/	0,
/* out0456_em-eta16-phi22*/	2,42,0,2,42,3,1,
/* out0457_em-eta17-phi22*/	1,42,0,6,
/* out0458_em-eta18-phi22*/	1,42,0,1,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	1,181,3,16,
/* out0461_em-eta1-phi23*/	1,181,2,15,
/* out0462_em-eta2-phi23*/	3,180,2,1,180,3,16,181,2,1,
/* out0463_em-eta3-phi23*/	6,112,0,4,112,2,2,113,0,12,113,1,2,179,3,2,180,2,15,
/* out0464_em-eta4-phi23*/	5,111,0,1,112,0,10,112,1,1,179,2,4,179,3,14,
/* out0465_em-eta5-phi23*/	3,111,0,10,178,5,5,179,2,12,
/* out0466_em-eta6-phi23*/	4,110,0,4,111,0,1,178,4,6,178,5,11,
/* out0467_em-eta7-phi23*/	3,110,0,4,178,3,7,178,4,10,
/* out0468_em-eta8-phi23*/	2,109,0,2,178,3,9,
/* out0469_em-eta9-phi23*/	1,109,0,1,
/* out0470_em-eta10-phi23*/	1,46,0,1,
/* out0471_em-eta11-phi23*/	1,46,0,3,
/* out0472_em-eta12-phi23*/	0,
/* out0473_em-eta13-phi23*/	0,
/* out0474_em-eta14-phi23*/	0,
/* out0475_em-eta15-phi23*/	0,
/* out0476_em-eta16-phi23*/	0,
/* out0477_em-eta17-phi23*/	0,
/* out0478_em-eta18-phi23*/	0,
/* out0479_em-eta19-phi23*/	0
};