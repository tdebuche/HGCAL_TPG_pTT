parameter integer matrixH [0:5849] = {
/* num inputs = 152(in0-in151) */
/* num outputs = 600(out0-out599) */
//* max inputs per outputs = 11 */
//* total number of input in adders 1749 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	0,
/* out0006_em-eta6-phi0*/	0,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	0,
/* out0010_em-eta10-phi0*/	0,
/* out0011_em-eta11-phi0*/	0,
/* out0012_em-eta12-phi0*/	0,
/* out0013_em-eta13-phi0*/	0,
/* out0014_em-eta14-phi0*/	0,
/* out0015_em-eta15-phi0*/	0,
/* out0016_em-eta16-phi0*/	0,
/* out0017_em-eta17-phi0*/	0,
/* out0018_em-eta18-phi0*/	0,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	0,
/* out0026_em-eta6-phi1*/	0,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	0,
/* out0029_em-eta9-phi1*/	0,
/* out0030_em-eta10-phi1*/	0,
/* out0031_em-eta11-phi1*/	0,
/* out0032_em-eta12-phi1*/	0,
/* out0033_em-eta13-phi1*/	0,
/* out0034_em-eta14-phi1*/	0,
/* out0035_em-eta15-phi1*/	0,
/* out0036_em-eta16-phi1*/	1,27,0,1,
/* out0037_em-eta17-phi1*/	0,
/* out0038_em-eta18-phi1*/	0,
/* out0039_em-eta19-phi1*/	1,12,5,2,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	0,
/* out0046_em-eta6-phi2*/	0,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	0,
/* out0049_em-eta9-phi2*/	0,
/* out0050_em-eta10-phi2*/	1,64,0,1,
/* out0051_em-eta11-phi2*/	0,
/* out0052_em-eta12-phi2*/	2,45,0,3,45,1,1,
/* out0053_em-eta13-phi2*/	2,45,0,12,45,3,2,
/* out0054_em-eta14-phi2*/	1,45,3,2,
/* out0055_em-eta15-phi2*/	2,27,0,2,27,1,7,
/* out0056_em-eta16-phi2*/	3,27,0,11,27,1,2,27,3,2,
/* out0057_em-eta17-phi2*/	2,27,0,2,27,3,9,
/* out0058_em-eta18-phi2*/	3,12,2,3,27,3,2,28,3,1,
/* out0059_em-eta19-phi2*/	3,12,2,5,12,4,1,12,5,9,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	2,119,1,2,119,2,3,
/* out0065_em-eta5-phi3*/	3,106,0,14,106,1,4,106,2,1,
/* out0066_em-eta6-phi3*/	4,93,0,7,93,1,4,106,0,2,106,2,3,
/* out0067_em-eta7-phi3*/	3,81,1,1,93,0,9,93,2,4,
/* out0068_em-eta8-phi3*/	2,81,0,11,81,1,3,
/* out0069_em-eta9-phi3*/	4,64,0,1,64,1,2,81,0,5,81,2,4,
/* out0070_em-eta10-phi3*/	2,64,0,9,64,1,2,
/* out0071_em-eta11-phi3*/	2,64,0,5,64,2,4,
/* out0072_em-eta12-phi3*/	4,45,1,13,45,2,2,46,0,3,46,1,12,
/* out0073_em-eta13-phi3*/	6,45,0,1,45,1,2,45,2,14,45,3,6,46,0,1,46,4,3,
/* out0074_em-eta14-phi3*/	4,28,1,3,45,3,6,46,3,12,46,4,1,
/* out0075_em-eta15-phi3*/	4,27,1,6,27,2,1,28,0,2,28,1,9,
/* out0076_em-eta16-phi3*/	4,27,1,1,27,2,12,28,0,2,28,4,1,
/* out0077_em-eta17-phi3*/	4,27,2,3,27,3,3,28,3,4,28,4,3,
/* out0078_em-eta18-phi3*/	3,12,2,5,12,3,1,28,3,7,
/* out0079_em-eta19-phi3*/	5,11,2,1,12,2,3,12,3,3,12,4,11,12,5,5,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	3,119,1,2,131,0,13,131,1,4,
/* out0084_em-eta4-phi4*/	6,119,1,12,119,2,13,120,0,8,120,1,2,131,0,3,131,2,2,
/* out0085_em-eta5-phi4*/	6,106,1,12,106,2,7,107,0,3,107,1,1,120,0,6,120,2,1,
/* out0086_em-eta6-phi4*/	3,93,1,10,106,2,5,107,0,9,
/* out0087_em-eta7-phi4*/	4,81,1,1,93,1,2,93,2,12,94,0,5,
/* out0088_em-eta8-phi4*/	3,81,1,11,81,2,3,94,0,2,
/* out0089_em-eta9-phi4*/	3,64,1,2,81,2,9,82,0,3,
/* out0090_em-eta10-phi4*/	2,64,1,9,64,2,2,
/* out0091_em-eta11-phi4*/	2,64,2,9,65,0,3,
/* out0092_em-eta12-phi4*/	5,45,4,15,45,5,6,46,0,5,46,1,4,65,0,2,
/* out0093_em-eta13-phi4*/	4,45,5,2,46,0,7,46,4,11,46,5,6,
/* out0094_em-eta14-phi4*/	5,27,4,3,46,2,14,46,3,4,46,4,1,46,5,1,
/* out0095_em-eta15-phi4*/	4,27,4,9,27,5,2,28,0,3,28,1,4,
/* out0096_em-eta16-phi4*/	3,27,5,1,28,0,9,28,4,6,
/* out0097_em-eta17-phi4*/	4,28,2,3,28,3,3,28,4,6,28,5,2,
/* out0098_em-eta18-phi4*/	3,12,3,6,28,2,6,28,3,1,
/* out0099_em-eta19-phi4*/	6,11,0,1,11,1,16,11,2,15,11,3,5,12,3,5,12,4,4,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	6,131,1,12,131,2,8,132,0,3,132,1,2,140,1,3,140,2,13,
/* out0104_em-eta4-phi5*/	6,120,0,1,120,1,14,120,2,3,121,0,1,131,2,6,132,0,11,
/* out0105_em-eta5-phi5*/	4,107,1,10,120,0,1,120,2,12,121,0,6,
/* out0106_em-eta6-phi5*/	4,107,0,4,107,1,5,107,2,15,108,0,1,
/* out0107_em-eta7-phi5*/	3,94,0,5,94,1,13,94,2,2,
/* out0108_em-eta8-phi5*/	4,82,0,1,82,1,4,94,0,4,94,2,8,
/* out0109_em-eta9-phi5*/	3,82,0,8,82,1,4,82,2,1,
/* out0110_em-eta10-phi5*/	6,64,1,1,64,2,1,65,1,2,66,1,7,82,0,4,82,2,4,
/* out0111_em-eta11-phi5*/	5,65,0,6,65,1,14,65,2,9,66,0,2,66,1,4,
/* out0112_em-eta12-phi5*/	6,45,4,1,45,5,4,65,0,5,65,2,4,65,3,15,66,3,3,
/* out0113_em-eta13-phi5*/	6,45,5,4,46,5,9,47,1,8,48,1,2,65,3,1,66,3,2,
/* out0114_em-eta14-phi5*/	5,46,2,2,47,0,12,47,1,6,47,2,1,47,3,1,
/* out0115_em-eta15-phi5*/	4,27,4,4,27,5,5,47,0,4,47,3,7,
/* out0116_em-eta16-phi5*/	2,27,5,8,28,5,7,
/* out0117_em-eta17-phi5*/	4,28,2,4,28,5,6,29,0,2,29,1,1,
/* out0118_em-eta18-phi5*/	4,11,3,2,12,3,1,28,2,3,29,0,6,
/* out0119_em-eta19-phi5*/	3,11,0,4,11,3,9,29,0,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	1,141,1,1,
/* out0123_em-eta3-phi6*/	6,132,1,11,140,1,13,140,2,3,141,0,16,141,1,3,141,2,1,
/* out0124_em-eta4-phi6*/	5,121,1,7,132,0,2,132,1,3,132,2,16,133,0,7,
/* out0125_em-eta5-phi6*/	3,121,0,9,121,1,8,121,2,13,
/* out0126_em-eta6-phi6*/	5,107,2,1,108,0,10,108,1,10,108,2,1,121,2,1,
/* out0127_em-eta7-phi6*/	6,94,1,3,94,2,3,95,0,2,95,1,3,108,0,5,108,2,5,
/* out0128_em-eta8-phi6*/	3,82,1,2,94,2,3,95,0,11,
/* out0129_em-eta9-phi6*/	4,82,1,6,82,2,6,83,0,1,95,0,1,
/* out0130_em-eta10-phi6*/	4,65,4,13,66,1,2,82,2,5,83,0,3,
/* out0131_em-eta11-phi6*/	7,65,2,2,65,4,3,65,5,9,66,0,14,66,1,3,66,4,6,66,5,2,
/* out0132_em-eta12-phi6*/	5,65,2,1,66,2,9,66,3,10,66,4,10,66,5,3,
/* out0133_em-eta13-phi6*/	5,47,1,1,47,4,5,48,0,4,48,1,14,66,3,1,
/* out0134_em-eta14-phi6*/	4,47,1,1,47,2,13,48,0,5,48,4,3,
/* out0135_em-eta15-phi6*/	4,47,2,2,47,3,7,48,3,7,48,4,3,
/* out0136_em-eta16-phi6*/	5,28,5,1,29,1,3,30,1,6,47,3,1,48,3,3,
/* out0137_em-eta17-phi6*/	3,29,1,11,29,2,2,30,1,1,
/* out0138_em-eta18-phi6*/	4,29,0,5,29,1,1,29,2,2,29,3,3,
/* out0139_em-eta19-phi6*/	3,11,0,11,29,0,2,29,3,7,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	4,141,1,3,148,0,9,148,1,3,148,2,6,
/* out0143_em-eta3-phi7*/	8,133,1,3,141,1,9,141,2,15,142,0,10,142,1,2,148,0,6,148,1,11,148,2,7,
/* out0144_em-eta4-phi7*/	4,133,0,8,133,1,13,133,2,13,142,0,1,
/* out0145_em-eta5-phi7*/	7,121,1,1,121,2,2,122,0,11,122,1,10,122,2,2,133,0,1,133,2,2,
/* out0146_em-eta6-phi7*/	6,108,1,6,108,2,5,109,0,3,109,1,2,122,0,5,122,2,3,
/* out0147_em-eta7-phi7*/	3,95,1,9,108,2,5,109,0,7,
/* out0148_em-eta8-phi7*/	3,95,0,2,95,1,4,95,2,11,
/* out0149_em-eta9-phi7*/	3,83,0,2,83,1,8,95,2,3,
/* out0150_em-eta10-phi7*/	3,83,0,9,83,1,1,83,2,2,
/* out0151_em-eta11-phi7*/	6,65,5,7,66,5,8,67,1,7,68,1,4,83,0,1,83,2,2,
/* out0152_em-eta12-phi7*/	6,47,4,1,66,2,7,66,5,3,67,0,13,67,1,8,67,3,1,
/* out0153_em-eta13-phi7*/	5,47,4,10,47,5,10,48,0,2,67,0,3,67,3,2,
/* out0154_em-eta14-phi7*/	4,47,5,2,48,0,5,48,4,8,48,5,7,
/* out0155_em-eta15-phi7*/	4,48,2,11,48,3,5,48,4,2,48,5,1,
/* out0156_em-eta16-phi7*/	3,29,4,6,30,1,8,48,3,1,
/* out0157_em-eta17-phi7*/	3,29,2,3,30,0,9,30,1,1,
/* out0158_em-eta18-phi7*/	3,29,2,8,29,3,1,30,4,3,
/* out0159_em-eta19-phi7*/	4,29,2,1,29,3,5,30,3,4,30,4,1,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	2,149,0,14,149,1,7,
/* out0163_em-eta3-phi8*/	11,142,0,4,142,1,14,142,2,12,143,0,2,143,2,5,148,0,1,148,1,2,148,2,3,149,0,2,149,1,1,149,2,12,
/* out0164_em-eta4-phi8*/	7,133,2,1,134,0,12,134,1,13,134,2,4,142,0,1,142,2,4,143,2,1,
/* out0165_em-eta5-phi8*/	6,122,1,6,122,2,7,123,0,5,123,1,3,134,0,4,134,2,4,
/* out0166_em-eta6-phi8*/	4,109,1,13,109,2,1,122,2,4,123,0,5,
/* out0167_em-eta7-phi8*/	3,96,1,2,109,0,6,109,2,12,
/* out0168_em-eta8-phi8*/	3,95,2,2,96,0,10,96,1,4,
/* out0169_em-eta9-phi8*/	3,83,1,7,83,2,1,96,0,6,
/* out0170_em-eta10-phi8*/	2,83,2,10,84,0,1,
/* out0171_em-eta11-phi8*/	5,67,4,12,67,5,1,68,0,7,68,1,12,83,2,1,
/* out0172_em-eta12-phi8*/	5,67,1,1,67,2,16,67,3,2,68,0,6,68,4,7,
/* out0173_em-eta13-phi8*/	5,47,5,3,50,1,2,67,3,11,68,3,10,68,4,1,
/* out0174_em-eta14-phi8*/	5,47,5,1,48,2,1,48,5,8,49,1,11,50,1,2,
/* out0175_em-eta15-phi8*/	4,29,4,1,48,2,4,49,0,12,49,1,2,
/* out0176_em-eta16-phi8*/	3,29,4,9,29,5,5,49,0,2,
/* out0177_em-eta17-phi8*/	3,29,5,3,30,0,7,30,4,3,
/* out0178_em-eta18-phi8*/	4,30,2,1,30,3,5,30,4,9,30,5,1,
/* out0179_em-eta19-phi8*/	2,30,2,2,30,3,7,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	1,149,1,5,
/* out0183_em-eta3-phi9*/	5,143,0,14,143,1,11,143,2,6,149,1,3,149,2,4,
/* out0184_em-eta4-phi9*/	6,134,1,3,134,2,6,135,0,9,135,1,8,143,1,5,143,2,4,
/* out0185_em-eta5-phi9*/	5,123,0,2,123,1,13,123,2,6,134,2,2,135,0,7,
/* out0186_em-eta6-phi9*/	6,109,1,1,109,2,1,110,0,1,110,1,7,123,0,4,123,2,10,
/* out0187_em-eta7-phi9*/	4,96,1,3,109,2,2,110,0,14,110,1,1,
/* out0188_em-eta8-phi9*/	3,96,1,7,96,2,9,110,0,1,
/* out0189_em-eta9-phi9*/	3,84,0,1,84,1,6,96,2,7,
/* out0190_em-eta10-phi9*/	2,84,0,10,84,1,2,
/* out0191_em-eta11-phi9*/	5,67,4,4,67,5,15,68,0,1,68,5,3,84,0,4,
/* out0192_em-eta12-phi9*/	5,68,0,2,68,2,8,68,3,1,68,4,8,68,5,13,
/* out0193_em-eta13-phi9*/	4,49,4,8,50,1,5,68,2,8,68,3,5,
/* out0194_em-eta14-phi9*/	4,49,1,2,49,2,5,50,0,8,50,1,7,
/* out0195_em-eta15-phi9*/	4,49,0,1,49,1,1,49,2,11,49,3,5,
/* out0196_em-eta16-phi9*/	3,29,5,4,49,0,1,49,3,11,
/* out0197_em-eta17-phi9*/	2,29,5,4,30,5,9,
/* out0198_em-eta18-phi9*/	2,30,2,5,30,5,6,
/* out0199_em-eta19-phi9*/	1,30,2,8,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	2,150,0,8,150,1,3,
/* out0203_em-eta3-phi10*/	5,144,0,15,144,1,11,144,2,3,150,0,8,150,2,5,
/* out0204_em-eta4-phi10*/	6,135,1,8,135,2,9,136,0,6,136,1,3,144,0,1,144,2,12,
/* out0205_em-eta5-phi10*/	5,124,0,6,124,1,13,124,2,1,135,2,7,136,0,2,
/* out0206_em-eta6-phi10*/	6,110,1,7,110,2,1,111,0,1,111,1,1,124,0,10,124,2,4,
/* out0207_em-eta7-phi10*/	4,97,1,3,110,1,1,110,2,14,111,0,2,
/* out0208_em-eta8-phi10*/	3,97,0,9,97,1,7,110,2,1,
/* out0209_em-eta9-phi10*/	3,84,1,6,84,2,1,97,0,7,
/* out0210_em-eta10-phi10*/	2,84,1,2,84,2,10,
/* out0211_em-eta11-phi10*/	5,69,1,3,69,4,4,70,0,1,70,1,15,84,2,4,
/* out0212_em-eta12-phi10*/	5,69,0,8,69,1,13,69,2,8,69,3,1,70,0,2,
/* out0213_em-eta13-phi10*/	4,49,4,8,49,5,5,69,0,8,69,3,5,
/* out0214_em-eta14-phi10*/	4,49,5,7,50,0,8,50,4,5,50,5,2,
/* out0215_em-eta15-phi10*/	4,50,2,1,50,3,5,50,4,11,50,5,1,
/* out0216_em-eta16-phi10*/	3,32,1,4,50,2,1,50,3,11,
/* out0217_em-eta17-phi10*/	2,31,1,9,32,1,4,
/* out0218_em-eta18-phi10*/	2,31,0,5,31,1,6,
/* out0219_em-eta19-phi10*/	1,31,0,8,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	1,150,1,11,
/* out0223_em-eta3-phi11*/	9,144,1,5,145,0,12,145,1,14,145,2,4,150,1,2,150,2,11,151,0,3,151,1,2,151,2,1,
/* out0224_em-eta4-phi11*/	7,136,0,4,136,1,13,136,2,12,137,0,1,144,2,1,145,0,4,145,2,1,
/* out0225_em-eta5-phi11*/	6,124,1,3,124,2,5,125,0,7,125,1,6,136,0,4,136,2,4,
/* out0226_em-eta6-phi11*/	4,111,0,1,111,1,13,124,2,6,125,0,4,
/* out0227_em-eta7-phi11*/	3,97,1,2,111,0,12,111,2,6,
/* out0228_em-eta8-phi11*/	3,97,1,4,97,2,10,98,0,2,
/* out0229_em-eta9-phi11*/	3,85,0,1,85,1,7,97,2,6,
/* out0230_em-eta10-phi11*/	2,84,2,1,85,0,10,
/* out0231_em-eta11-phi11*/	5,69,4,12,69,5,12,70,0,7,70,1,1,85,0,1,
/* out0232_em-eta12-phi11*/	5,69,2,7,70,0,6,70,3,2,70,4,16,70,5,1,
/* out0233_em-eta13-phi11*/	5,49,5,2,52,1,3,69,2,1,69,3,10,70,3,11,
/* out0234_em-eta14-phi11*/	5,49,5,2,50,5,11,51,0,1,51,1,8,52,1,1,
/* out0235_em-eta15-phi11*/	4,31,4,1,50,2,12,50,5,2,51,0,4,
/* out0236_em-eta16-phi11*/	3,31,4,9,32,1,5,50,2,2,
/* out0237_em-eta17-phi11*/	3,31,2,3,32,0,7,32,1,3,
/* out0238_em-eta18-phi11*/	4,31,0,1,31,1,1,31,2,9,31,3,5,
/* out0239_em-eta19-phi11*/	2,31,0,2,31,3,7,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	4,146,1,3,151,0,6,151,1,3,151,2,9,
/* out0243_em-eta3-phi12*/	8,137,1,3,145,1,2,145,2,10,146,0,15,146,1,9,151,0,7,151,1,11,151,2,6,
/* out0244_em-eta4-phi12*/	4,137,0,13,137,1,13,137,2,8,145,2,1,
/* out0245_em-eta5-phi12*/	7,125,0,2,125,1,10,125,2,11,126,0,2,126,1,1,137,0,2,137,2,1,
/* out0246_em-eta6-phi12*/	6,111,1,2,111,2,3,112,0,5,112,1,6,125,0,3,125,2,5,
/* out0247_em-eta7-phi12*/	3,98,1,9,111,2,7,112,0,5,
/* out0248_em-eta8-phi12*/	3,98,0,11,98,1,4,98,2,2,
/* out0249_em-eta9-phi12*/	3,85,1,8,85,2,2,98,0,3,
/* out0250_em-eta10-phi12*/	3,85,0,2,85,1,1,85,2,9,
/* out0251_em-eta11-phi12*/	6,69,5,4,70,5,7,71,1,8,72,1,7,85,0,2,85,2,1,
/* out0252_em-eta12-phi12*/	6,51,4,1,70,2,13,70,3,1,70,5,8,71,0,7,71,1,3,
/* out0253_em-eta13-phi12*/	5,51,4,10,52,0,2,52,1,10,70,2,3,70,3,2,
/* out0254_em-eta14-phi12*/	4,51,1,7,51,2,8,52,0,5,52,1,2,
/* out0255_em-eta15-phi12*/	4,51,0,11,51,1,1,51,2,2,51,3,5,
/* out0256_em-eta16-phi12*/	3,31,4,6,31,5,8,51,3,1,
/* out0257_em-eta17-phi12*/	3,31,5,1,32,0,9,32,4,3,
/* out0258_em-eta18-phi12*/	3,31,2,3,32,3,1,32,4,8,
/* out0259_em-eta19-phi12*/	4,31,2,1,31,3,4,32,3,5,32,4,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	1,146,1,1,
/* out0263_em-eta3-phi13*/	6,138,1,11,146,0,1,146,1,3,146,2,16,147,0,12,147,2,4,
/* out0264_em-eta4-phi13*/	5,126,1,7,137,2,7,138,0,16,138,1,3,138,2,2,
/* out0265_em-eta5-phi13*/	3,126,0,13,126,1,8,126,2,9,
/* out0266_em-eta6-phi13*/	5,112,0,1,112,1,10,112,2,10,113,0,1,126,0,1,
/* out0267_em-eta7-phi13*/	6,98,1,3,98,2,2,99,0,3,99,1,3,112,0,5,112,2,5,
/* out0268_em-eta8-phi13*/	3,86,1,2,98,2,11,99,0,3,
/* out0269_em-eta9-phi13*/	4,85,2,1,86,0,6,86,1,6,98,2,1,
/* out0270_em-eta10-phi13*/	4,71,4,13,71,5,2,85,2,3,86,0,5,
/* out0271_em-eta11-phi13*/	7,71,1,2,71,2,6,71,4,3,71,5,3,72,0,14,72,1,9,72,4,2,
/* out0272_em-eta12-phi13*/	5,71,0,9,71,1,3,71,2,10,71,3,10,72,4,1,
/* out0273_em-eta13-phi13*/	5,51,4,5,51,5,14,52,0,4,52,5,1,71,3,1,
/* out0274_em-eta14-phi13*/	4,51,2,3,52,0,5,52,4,13,52,5,1,
/* out0275_em-eta15-phi13*/	4,51,2,3,51,3,7,52,3,7,52,4,2,
/* out0276_em-eta16-phi13*/	5,31,5,6,32,5,3,33,1,1,51,3,3,52,3,1,
/* out0277_em-eta17-phi13*/	3,31,5,1,32,4,2,32,5,11,
/* out0278_em-eta18-phi13*/	4,32,2,5,32,3,3,32,4,2,32,5,1,
/* out0279_em-eta19-phi13*/	3,13,4,11,32,2,2,32,3,7,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	6,138,1,2,138,2,3,139,0,8,139,1,12,147,0,4,147,2,12,
/* out0284_em-eta4-phi14*/	6,126,2,1,127,0,3,127,1,14,127,2,1,138,2,11,139,0,6,
/* out0285_em-eta5-phi14*/	4,113,1,10,126,2,6,127,0,12,127,2,1,
/* out0286_em-eta6-phi14*/	4,112,2,1,113,0,15,113,1,5,113,2,4,
/* out0287_em-eta7-phi14*/	3,99,0,2,99,1,13,99,2,5,
/* out0288_em-eta8-phi14*/	4,86,1,4,86,2,1,99,0,8,99,2,4,
/* out0289_em-eta9-phi14*/	3,86,0,1,86,1,4,86,2,8,
/* out0290_em-eta10-phi14*/	6,71,5,7,72,5,2,73,0,1,73,1,1,86,0,4,86,2,4,
/* out0291_em-eta11-phi14*/	5,71,5,4,72,0,2,72,2,6,72,4,9,72,5,14,
/* out0292_em-eta12-phi14*/	6,53,4,1,54,1,4,71,3,3,72,2,5,72,3,15,72,4,4,
/* out0293_em-eta13-phi14*/	6,51,5,2,52,5,8,53,1,9,54,1,4,71,3,2,72,3,1,
/* out0294_em-eta14-phi14*/	5,52,2,12,52,3,1,52,4,1,52,5,6,53,0,2,
/* out0295_em-eta15-phi14*/	4,33,4,4,34,1,5,52,2,4,52,3,7,
/* out0296_em-eta16-phi14*/	2,33,1,7,34,1,8,
/* out0297_em-eta17-phi14*/	4,32,2,2,32,5,1,33,0,4,33,1,6,
/* out0298_em-eta18-phi14*/	4,13,5,2,14,5,1,32,2,6,33,0,3,
/* out0299_em-eta19-phi14*/	3,13,4,4,13,5,9,32,2,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	2,139,1,4,139,2,13,
/* out0304_em-eta4-phi15*/	5,127,1,2,127,2,8,128,2,5,139,0,2,139,2,3,
/* out0305_em-eta5-phi15*/	6,113,1,1,113,2,3,114,0,7,114,1,12,127,0,1,127,2,6,
/* out0306_em-eta6-phi15*/	3,100,1,10,113,2,9,114,0,5,
/* out0307_em-eta7-phi15*/	4,87,1,1,99,2,5,100,0,12,100,1,2,
/* out0308_em-eta8-phi15*/	3,87,0,3,87,1,11,99,2,2,
/* out0309_em-eta9-phi15*/	3,73,1,2,86,2,3,87,0,9,
/* out0310_em-eta10-phi15*/	2,73,0,2,73,1,9,
/* out0311_em-eta11-phi15*/	2,72,2,3,73,0,9,
/* out0312_em-eta12-phi15*/	5,53,4,15,53,5,4,54,0,5,54,1,6,72,2,2,
/* out0313_em-eta13-phi15*/	4,53,1,6,53,2,11,54,0,7,54,1,2,
/* out0314_em-eta14-phi15*/	5,33,4,3,53,0,14,53,1,1,53,2,1,53,3,4,
/* out0315_em-eta15-phi15*/	4,33,4,9,33,5,4,34,0,3,34,1,2,
/* out0316_em-eta16-phi15*/	3,33,2,6,34,0,9,34,1,1,
/* out0317_em-eta17-phi15*/	4,33,0,3,33,1,2,33,2,6,33,3,3,
/* out0318_em-eta18-phi15*/	3,14,5,6,33,0,6,33,3,1,
/* out0319_em-eta19-phi15*/	6,13,4,1,13,5,5,14,0,15,14,1,16,14,4,4,14,5,5,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	4,128,1,1,128,2,1,129,0,6,129,1,12,
/* out0324_em-eta4-phi16*/	5,115,0,1,115,1,9,128,1,15,128,2,10,129,0,5,
/* out0325_em-eta5-phi16*/	5,101,1,3,114,0,1,114,1,4,114,2,14,115,0,7,
/* out0326_em-eta6-phi16*/	6,100,1,4,100,2,7,101,0,6,101,1,4,114,0,3,114,2,2,
/* out0327_em-eta7-phi16*/	5,87,1,1,88,0,1,88,1,4,100,0,4,100,2,9,
/* out0328_em-eta8-phi16*/	3,87,1,3,87,2,11,88,0,2,
/* out0329_em-eta9-phi16*/	6,73,1,2,73,2,1,74,0,1,74,1,2,87,0,4,87,2,5,
/* out0330_em-eta10-phi16*/	2,73,1,2,73,2,9,
/* out0331_em-eta11-phi16*/	3,56,1,3,73,0,4,73,2,5,
/* out0332_em-eta12-phi16*/	5,53,5,12,54,0,3,54,4,2,54,5,13,55,1,2,
/* out0333_em-eta13-phi16*/	6,53,2,3,54,0,1,54,2,1,54,3,6,54,4,14,54,5,2,
/* out0334_em-eta14-phi16*/	4,33,5,3,53,2,1,53,3,12,54,3,6,
/* out0335_em-eta15-phi16*/	4,33,5,9,34,0,2,34,4,1,34,5,6,
/* out0336_em-eta16-phi16*/	4,33,2,1,34,0,2,34,4,12,34,5,1,
/* out0337_em-eta17-phi16*/	4,33,2,3,33,3,4,34,3,3,34,4,3,
/* out0338_em-eta18-phi16*/	3,14,2,5,14,5,1,33,3,7,
/* out0339_em-eta19-phi16*/	5,14,0,1,14,2,3,14,3,5,14,4,11,14,5,3,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	6,116,1,5,129,0,1,129,1,4,129,2,14,130,0,13,130,2,3,
/* out0344_em-eta4-phi17*/	6,115,1,7,115,2,11,116,0,7,116,1,4,129,0,4,129,2,2,
/* out0345_em-eta5-phi17*/	6,101,1,6,101,2,4,102,0,3,102,1,4,115,0,8,115,2,5,
/* out0346_em-eta6-phi17*/	3,101,0,10,101,1,3,101,2,10,
/* out0347_em-eta7-phi17*/	3,88,0,2,88,1,12,88,2,6,
/* out0348_em-eta8-phi17*/	3,74,1,4,88,0,11,88,2,1,
/* out0349_em-eta9-phi17*/	3,74,0,4,74,1,9,74,2,1,
/* out0350_em-eta10-phi17*/	4,55,4,8,55,5,2,73,2,1,74,0,8,
/* out0351_em-eta11-phi17*/	6,55,1,1,55,2,2,55,4,8,55,5,2,56,0,9,56,1,13,
/* out0352_em-eta12-phi17*/	5,54,2,3,54,5,1,55,0,10,55,1,13,55,2,5,
/* out0353_em-eta13-phi17*/	5,35,4,10,36,1,1,54,2,12,54,3,2,55,0,3,
/* out0354_em-eta14-phi17*/	3,35,1,5,36,1,14,54,3,2,
/* out0355_em-eta15-phi17*/	4,34,2,2,34,5,7,35,0,3,35,1,8,
/* out0356_em-eta16-phi17*/	3,34,2,11,34,3,2,34,5,2,
/* out0357_em-eta17-phi17*/	4,15,4,1,16,1,2,34,2,2,34,3,9,
/* out0358_em-eta18-phi17*/	5,14,2,3,15,1,3,16,1,4,33,3,1,34,3,2,
/* out0359_em-eta19-phi17*/	4,14,2,5,14,3,9,14,4,1,15,1,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	1,117,1,2,
/* out0363_em-eta3-phi18*/	6,116,1,5,116,2,6,117,0,9,117,1,11,130,0,3,130,2,13,
/* out0364_em-eta4-phi18*/	7,102,1,5,102,2,2,103,0,2,103,1,5,116,0,9,116,1,2,116,2,10,
/* out0365_em-eta5-phi18*/	3,102,0,12,102,1,7,102,2,11,
/* out0366_em-eta6-phi18*/	5,89,0,3,89,1,16,89,2,3,101,2,2,102,0,1,
/* out0367_em-eta7-phi18*/	3,75,1,4,88,2,6,89,0,10,
/* out0368_em-eta8-phi18*/	5,74,1,1,74,2,2,75,0,5,75,1,6,88,2,3,
/* out0369_em-eta9-phi18*/	3,57,1,1,74,2,11,75,0,2,
/* out0370_em-eta10-phi18*/	6,55,5,9,56,5,6,57,0,1,57,1,2,74,0,3,74,2,2,
/* out0371_em-eta11-phi18*/	7,55,2,2,55,5,3,56,0,7,56,2,1,56,3,2,56,4,14,56,5,10,
/* out0372_em-eta12-phi18*/	5,55,0,2,55,2,7,55,3,15,56,3,5,56,4,2,
/* out0373_em-eta13-phi18*/	4,35,4,6,35,5,13,36,0,5,55,0,1,
/* out0374_em-eta14-phi18*/	4,35,2,8,36,0,11,36,1,1,36,4,2,
/* out0375_em-eta15-phi18*/	4,35,0,8,35,1,3,35,2,5,35,3,3,
/* out0376_em-eta16-phi18*/	3,15,4,10,34,2,1,35,0,5,
/* out0377_em-eta17-phi18*/	3,15,4,4,16,0,2,16,1,7,
/* out0378_em-eta18-phi18*/	4,15,1,5,15,2,1,16,0,1,16,1,3,
/* out0379_em-eta19-phi18*/	3,14,3,2,15,0,3,15,1,5,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	5,117,1,1,117,2,1,118,0,9,118,1,3,118,2,6,
/* out0383_em-eta3-phi19*/	10,103,1,2,103,2,1,104,0,3,104,1,9,117,0,7,117,1,2,117,2,15,118,0,6,118,1,11,118,2,7,
/* out0384_em-eta4-phi19*/	4,103,0,11,103,1,9,103,2,14,104,0,1,
/* out0385_em-eta5-phi19*/	5,90,0,5,90,1,16,90,2,3,102,2,3,103,0,3,
/* out0386_em-eta6-phi19*/	3,76,1,5,89,2,11,90,0,8,
/* out0387_em-eta7-phi19*/	6,75,1,4,75,2,5,76,0,4,76,1,3,89,0,3,89,2,2,
/* out0388_em-eta8-phi19*/	3,75,0,6,75,1,2,75,2,9,
/* out0389_em-eta9-phi19*/	3,57,1,10,57,2,1,75,0,3,
/* out0390_em-eta10-phi19*/	2,57,0,8,57,1,3,
/* out0391_em-eta11-phi19*/	4,37,4,11,56,2,14,56,3,1,57,0,3,
/* out0392_em-eta12-phi19*/	7,35,5,1,37,1,5,37,4,1,38,1,15,55,3,1,56,2,1,56,3,8,
/* out0393_em-eta13-phi19*/	6,35,5,2,36,2,3,36,4,2,36,5,15,37,0,1,37,1,5,
/* out0394_em-eta14-phi19*/	5,35,2,1,36,2,3,36,3,6,36,4,12,36,5,1,
/* out0395_em-eta15-phi19*/	3,35,2,2,35,3,12,36,3,4,
/* out0396_em-eta16-phi19*/	3,15,4,1,15,5,13,35,3,1,
/* out0397_em-eta17-phi19*/	3,15,5,1,16,0,11,16,4,1,
/* out0398_em-eta18-phi19*/	2,15,2,9,16,0,2,
/* out0399_em-eta19-phi19*/	4,15,0,5,15,1,2,15,2,2,15,3,1,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	1,105,1,12,
/* out0403_em-eta3-phi20*/	11,92,0,2,92,2,5,104,0,7,104,1,7,104,2,16,105,0,16,105,1,1,105,2,5,118,0,1,118,1,2,118,2,3,
/* out0404_em-eta4-phi20*/	6,91,0,6,91,1,16,91,2,7,92,2,1,103,2,1,104,0,5,
/* out0405_em-eta5-phi20*/	3,77,1,8,90,2,12,91,0,9,
/* out0406_em-eta6-phi20*/	6,76,1,7,76,2,8,77,0,4,77,1,2,90,0,3,90,2,1,
/* out0407_em-eta7-phi20*/	4,58,1,2,76,0,12,76,1,1,76,2,4,
/* out0408_em-eta8-phi20*/	3,58,0,2,58,1,12,75,2,2,
/* out0409_em-eta9-phi20*/	2,57,2,8,58,0,6,
/* out0410_em-eta10-phi20*/	3,39,1,1,57,0,3,57,2,7,
/* out0411_em-eta11-phi20*/	6,37,4,4,37,5,16,38,0,5,38,4,2,38,5,6,57,0,1,
/* out0412_em-eta12-phi20*/	5,37,1,2,37,2,13,38,0,11,38,1,1,38,4,5,
/* out0413_em-eta13-phi20*/	6,17,4,2,36,2,3,37,0,14,37,1,4,37,2,1,37,3,3,
/* out0414_em-eta14-phi20*/	4,17,4,9,18,1,4,36,2,7,36,3,2,
/* out0415_em-eta15-phi20*/	4,16,5,1,17,1,4,18,1,9,36,3,4,
/* out0416_em-eta16-phi20*/	3,15,5,2,16,5,12,17,1,2,
/* out0417_em-eta17-phi20*/	2,16,4,10,16,5,3,
/* out0418_em-eta18-phi20*/	4,15,2,4,15,3,1,16,3,1,16,4,5,
/* out0419_em-eta19-phi20*/	2,15,0,8,15,3,9,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	2,105,1,3,105,2,4,
/* out0423_em-eta3-phi21*/	4,92,0,14,92,1,11,92,2,6,105,2,7,
/* out0424_em-eta4-phi21*/	5,78,0,2,78,1,16,91,2,8,92,1,5,92,2,4,
/* out0425_em-eta5-phi21*/	5,77,1,6,77,2,14,78,0,6,91,0,1,91,2,1,
/* out0426_em-eta6-phi21*/	4,59,1,9,76,2,2,77,0,12,77,2,2,
/* out0427_em-eta7-phi21*/	5,58,1,1,58,2,2,59,0,8,59,1,7,76,2,2,
/* out0428_em-eta8-phi21*/	3,58,0,2,58,1,1,58,2,13,
/* out0429_em-eta9-phi21*/	3,39,1,7,58,0,6,58,2,1,
/* out0430_em-eta10-phi21*/	2,39,0,4,39,1,8,
/* out0431_em-eta11-phi21*/	4,38,2,11,38,4,1,38,5,10,39,0,4,
/* out0432_em-eta12-phi21*/	5,37,2,2,37,3,2,38,2,5,38,3,15,38,4,8,
/* out0433_em-eta13-phi21*/	5,17,4,2,17,5,11,37,0,1,37,3,11,38,3,1,
/* out0434_em-eta14-phi21*/	4,17,4,3,17,5,5,18,0,13,18,1,2,
/* out0435_em-eta15-phi21*/	4,17,1,6,17,2,8,18,0,3,18,1,1,
/* out0436_em-eta16-phi21*/	3,16,2,4,17,0,8,17,1,4,
/* out0437_em-eta17-phi21*/	2,16,2,12,16,3,2,
/* out0438_em-eta18-phi21*/	1,16,3,10,
/* out0439_em-eta19-phi21*/	2,15,3,5,16,3,3,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	1,80,1,7,
/* out0443_em-eta3-phi22*/	5,79,0,3,79,1,15,79,2,5,80,0,11,80,1,3,
/* out0444_em-eta4-phi22*/	5,61,1,8,78,0,2,78,2,16,79,0,13,79,2,5,
/* out0445_em-eta5-phi22*/	5,60,1,14,60,2,6,61,0,1,61,1,1,78,0,6,
/* out0446_em-eta6-phi22*/	4,41,1,2,59,2,9,60,0,12,60,1,2,
/* out0447_em-eta7-phi22*/	5,40,1,2,40,2,1,41,1,2,59,0,8,59,2,7,
/* out0448_em-eta8-phi22*/	3,40,0,2,40,1,13,40,2,1,
/* out0449_em-eta9-phi22*/	3,39,2,7,40,0,6,40,1,1,
/* out0450_em-eta10-phi22*/	2,39,0,4,39,2,8,
/* out0451_em-eta11-phi22*/	4,19,4,11,19,5,10,20,0,1,39,0,4,
/* out0452_em-eta12-phi22*/	5,19,1,2,19,2,2,19,4,5,20,0,8,20,1,15,
/* out0453_em-eta13-phi22*/	5,18,2,2,18,5,11,19,0,1,19,1,11,20,1,1,
/* out0454_em-eta14-phi22*/	4,18,2,3,18,3,2,18,4,13,18,5,5,
/* out0455_em-eta15-phi22*/	4,17,2,8,17,3,6,18,3,1,18,4,3,
/* out0456_em-eta16-phi22*/	3,0,4,4,17,0,8,17,3,4,
/* out0457_em-eta17-phi22*/	2,0,4,12,1,1,2,
/* out0458_em-eta18-phi22*/	1,1,1,10,
/* out0459_em-eta19-phi22*/	2,0,1,5,1,1,3,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	2,80,1,6,80,2,6,
/* out0463_em-eta3-phi23*/	10,62,0,7,62,1,16,62,2,7,63,0,3,63,1,2,63,2,1,79,1,1,79,2,5,80,0,5,80,2,10,
/* out0464_em-eta4-phi23*/	6,43,1,1,61,0,6,61,1,7,61,2,16,62,0,5,79,2,1,
/* out0465_em-eta5-phi23*/	3,42,1,12,60,2,8,61,0,9,
/* out0466_em-eta6-phi23*/	6,41,1,8,41,2,7,42,0,3,42,1,1,60,0,4,60,2,2,
/* out0467_em-eta7-phi23*/	4,40,2,2,41,0,12,41,1,4,41,2,1,
/* out0468_em-eta8-phi23*/	3,22,1,2,40,0,2,40,2,12,
/* out0469_em-eta9-phi23*/	2,21,1,8,40,0,6,
/* out0470_em-eta10-phi23*/	3,21,0,3,21,1,7,39,2,1,
/* out0471_em-eta11-phi23*/	6,19,5,6,20,0,2,20,2,4,20,4,5,20,5,16,21,0,1,
/* out0472_em-eta12-phi23*/	5,19,2,13,19,3,2,20,0,5,20,3,1,20,4,11,
/* out0473_em-eta13-phi23*/	6,2,4,3,18,2,2,19,0,14,19,1,3,19,2,1,19,3,4,
/* out0474_em-eta14-phi23*/	4,2,4,7,3,1,2,18,2,9,18,3,4,
/* out0475_em-eta15-phi23*/	4,0,5,1,3,1,4,17,3,4,18,3,9,
/* out0476_em-eta16-phi23*/	3,0,5,12,1,5,2,17,3,2,
/* out0477_em-eta17-phi23*/	2,0,5,3,1,0,10,
/* out0478_em-eta18-phi23*/	4,0,1,1,0,2,4,1,0,5,1,1,1,
/* out0479_em-eta19-phi23*/	2,0,0,8,0,1,9,
/* out0480_em-eta0-phi24*/	0,
/* out0481_em-eta1-phi24*/	0,
/* out0482_em-eta2-phi24*/	5,44,1,1,44,2,1,63,0,6,63,1,3,63,2,9,
/* out0483_em-eta3-phi24*/	10,43,1,1,43,2,2,44,0,7,44,1,15,44,2,2,62,0,3,62,2,9,63,0,7,63,1,11,63,2,6,
/* out0484_em-eta4-phi24*/	4,43,0,11,43,1,14,43,2,9,62,0,1,
/* out0485_em-eta5-phi24*/	5,24,1,3,42,0,5,42,1,3,42,2,16,43,0,3,
/* out0486_em-eta6-phi24*/	3,23,1,11,41,2,5,42,0,8,
/* out0487_em-eta7-phi24*/	6,22,1,5,22,2,4,23,0,3,23,1,2,41,0,4,41,2,3,
/* out0488_em-eta8-phi24*/	3,22,0,6,22,1,9,22,2,2,
/* out0489_em-eta9-phi24*/	3,21,1,1,21,2,10,22,0,3,
/* out0490_em-eta10-phi24*/	2,21,0,8,21,2,3,
/* out0491_em-eta11-phi24*/	4,4,4,14,5,1,1,20,2,11,21,0,3,
/* out0492_em-eta12-phi24*/	7,3,5,1,4,1,1,4,4,1,5,1,8,19,3,5,20,2,1,20,3,15,
/* out0493_em-eta13-phi24*/	6,2,4,3,2,5,15,3,0,2,3,5,2,19,0,1,19,3,5,
/* out0494_em-eta14-phi24*/	5,2,2,1,2,4,3,2,5,1,3,0,12,3,1,6,
/* out0495_em-eta15-phi24*/	3,2,1,12,2,2,2,3,1,4,
/* out0496_em-eta16-phi24*/	3,1,2,1,1,5,13,2,1,1,
/* out0497_em-eta17-phi24*/	3,1,0,1,1,4,11,1,5,1,
/* out0498_em-eta18-phi24*/	2,0,2,9,1,4,2,
/* out0499_em-eta19-phi24*/	4,0,0,5,0,1,1,0,2,2,0,3,2,
/* out0500_em-eta0-phi25*/	0,
/* out0501_em-eta1-phi25*/	0,
/* out0502_em-eta2-phi25*/	1,44,2,2,
/* out0503_em-eta3-phi25*/	6,25,1,6,25,2,5,26,0,12,26,2,4,44,0,9,44,2,11,
/* out0504_em-eta4-phi25*/	7,24,1,2,24,2,5,25,0,9,25,1,10,25,2,2,43,0,2,43,2,5,
/* out0505_em-eta5-phi25*/	3,24,0,12,24,1,11,24,2,7,
/* out0506_em-eta6-phi25*/	5,8,1,2,23,0,3,23,1,3,23,2,16,24,0,1,
/* out0507_em-eta7-phi25*/	3,7,1,6,22,2,4,23,0,10,
/* out0508_em-eta8-phi25*/	5,6,1,2,6,2,1,7,1,3,22,0,5,22,2,6,
/* out0509_em-eta9-phi25*/	3,6,1,11,21,2,1,22,0,2,
/* out0510_em-eta10-phi25*/	6,4,5,6,5,5,9,6,0,3,6,1,2,21,0,1,21,2,2,
/* out0511_em-eta11-phi25*/	7,4,2,2,4,4,1,4,5,10,5,0,14,5,1,2,5,4,7,5,5,3,
/* out0512_em-eta12-phi25*/	5,4,0,2,4,1,15,4,2,7,5,0,2,5,1,5,
/* out0513_em-eta13-phi25*/	4,3,2,6,3,4,5,3,5,13,4,0,1,
/* out0514_em-eta14-phi25*/	4,2,2,8,3,0,2,3,3,1,3,4,11,
/* out0515_em-eta15-phi25*/	4,2,0,8,2,1,3,2,2,5,2,3,3,
/* out0516_em-eta16-phi25*/	2,1,2,10,2,0,5,
/* out0517_em-eta17-phi25*/	3,1,2,4,1,3,7,1,4,2,
/* out0518_em-eta18-phi25*/	4,0,2,1,0,3,5,1,3,3,1,4,1,
/* out0519_em-eta19-phi25*/	2,0,0,3,0,3,5,
/* out0520_em-eta0-phi26*/	0,
/* out0521_em-eta1-phi26*/	0,
/* out0522_em-eta2-phi26*/	0,
/* out0523_em-eta3-phi26*/	6,10,0,1,10,1,14,10,2,4,25,2,5,26,0,4,26,2,12,
/* out0524_em-eta4-phi26*/	6,9,1,11,9,2,7,10,0,4,10,1,2,25,0,7,25,2,4,
/* out0525_em-eta5-phi26*/	6,8,1,4,8,2,6,9,0,8,9,1,5,24,0,3,24,2,4,
/* out0526_em-eta6-phi26*/	3,8,0,10,8,1,10,8,2,3,
/* out0527_em-eta7-phi26*/	3,7,0,2,7,1,6,7,2,12,
/* out0528_em-eta8-phi26*/	3,6,2,4,7,0,11,7,1,1,
/* out0529_em-eta9-phi26*/	3,6,0,4,6,1,1,6,2,9,
/* out0530_em-eta10-phi26*/	3,5,2,8,5,5,2,6,0,8,
/* out0531_em-eta11-phi26*/	6,4,2,2,4,3,1,5,2,8,5,3,13,5,4,9,5,5,2,
/* out0532_em-eta12-phi26*/	3,4,0,10,4,2,5,4,3,13,
/* out0533_em-eta13-phi26*/	3,3,2,10,3,3,1,4,0,3,
/* out0534_em-eta14-phi26*/	2,2,3,5,3,3,14,
/* out0535_em-eta15-phi26*/	2,2,0,3,2,3,8,
/* out0536_em-eta16-phi26*/	0,
/* out0537_em-eta17-phi26*/	2,1,2,1,1,3,2,
/* out0538_em-eta18-phi26*/	2,0,3,3,1,3,4,
/* out0539_em-eta19-phi26*/	1,0,3,1,
/* out0540_em-eta0-phi27*/	0,
/* out0541_em-eta1-phi27*/	0,
/* out0542_em-eta2-phi27*/	0,
/* out0543_em-eta3-phi27*/	2,10,0,6,10,2,12,
/* out0544_em-eta4-phi27*/	3,9,0,1,9,2,9,10,0,5,
/* out0545_em-eta5-phi27*/	2,8,2,3,9,0,7,
/* out0546_em-eta6-phi27*/	2,8,0,6,8,2,4,
/* out0547_em-eta7-phi27*/	2,7,0,1,7,2,4,
/* out0548_em-eta8-phi27*/	1,7,0,2,
/* out0549_em-eta9-phi27*/	2,6,0,1,6,2,2,
/* out0550_em-eta10-phi27*/	0,
/* out0551_em-eta11-phi27*/	1,5,3,3,
/* out0552_em-eta12-phi27*/	1,4,3,2,
/* out0553_em-eta13-phi27*/	0,
/* out0554_em-eta14-phi27*/	0,
/* out0555_em-eta15-phi27*/	0,
/* out0556_em-eta16-phi27*/	0,
/* out0557_em-eta17-phi27*/	0,
/* out0558_em-eta18-phi27*/	0,
/* out0559_em-eta19-phi27*/	0,
/* out0560_em-eta0-phi28*/	0,
/* out0561_em-eta1-phi28*/	0,
/* out0562_em-eta2-phi28*/	0,
/* out0563_em-eta3-phi28*/	0,
/* out0564_em-eta4-phi28*/	0,
/* out0565_em-eta5-phi28*/	0,
/* out0566_em-eta6-phi28*/	0,
/* out0567_em-eta7-phi28*/	0,
/* out0568_em-eta8-phi28*/	0,
/* out0569_em-eta9-phi28*/	0,
/* out0570_em-eta10-phi28*/	0,
/* out0571_em-eta11-phi28*/	0,
/* out0572_em-eta12-phi28*/	0,
/* out0573_em-eta13-phi28*/	0,
/* out0574_em-eta14-phi28*/	0,
/* out0575_em-eta15-phi28*/	0,
/* out0576_em-eta16-phi28*/	0,
/* out0577_em-eta17-phi28*/	0,
/* out0578_em-eta18-phi28*/	0,
/* out0579_em-eta19-phi28*/	0,
/* out0580_em-eta0-phi29*/	0,
/* out0581_em-eta1-phi29*/	0,
/* out0582_em-eta2-phi29*/	0,
/* out0583_em-eta3-phi29*/	0,
/* out0584_em-eta4-phi29*/	0,
/* out0585_em-eta5-phi29*/	0,
/* out0586_em-eta6-phi29*/	0,
/* out0587_em-eta7-phi29*/	0,
/* out0588_em-eta8-phi29*/	0,
/* out0589_em-eta9-phi29*/	0,
/* out0590_em-eta10-phi29*/	0,
/* out0591_em-eta11-phi29*/	0,
/* out0592_em-eta12-phi29*/	0,
/* out0593_em-eta13-phi29*/	0,
/* out0594_em-eta14-phi29*/	0,
/* out0595_em-eta15-phi29*/	0,
/* out0596_em-eta16-phi29*/	0,
/* out0597_em-eta17-phi29*/	0,
/* out0598_em-eta18-phi29*/	0,
/* out0599_em-eta19-phi29*/	0
};