parameter integer matrixH [0:10874] = {
/* num inputs = 322(in0-in321) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 14 */
//* total number of input in adders 3464 */

/* out0000_em-eta0-phi0*/	1,277,0,4,
/* out0001_em-eta1-phi0*/	2,277,0,12,277,1,6,
/* out0002_em-eta2-phi0*/	4,63,0,8,63,1,6,276,0,7,277,1,10,
/* out0003_em-eta3-phi0*/	6,62,0,7,62,1,4,63,0,8,63,2,5,276,0,9,276,1,9,
/* out0004_em-eta4-phi0*/	9,52,0,16,52,1,16,52,2,12,61,0,3,61,1,2,62,0,9,62,2,2,275,0,10,276,1,7,
/* out0005_em-eta5-phi0*/	8,51,0,16,51,1,16,51,2,6,52,2,4,61,0,11,61,2,1,275,0,6,275,1,11,
/* out0006_em-eta6-phi0*/	5,50,1,6,51,2,10,60,0,10,274,0,12,275,1,5,
/* out0007_em-eta7-phi0*/	7,50,0,16,50,1,10,50,2,14,59,0,3,60,0,1,274,0,4,274,1,13,
/* out0008_em-eta8-phi0*/	8,49,1,12,50,2,2,59,0,4,217,0,1,217,1,7,269,2,5,274,1,3,274,2,13,
/* out0009_em-eta9-phi0*/	13,48,1,2,49,0,16,49,1,1,49,2,12,58,0,2,217,0,7,217,1,5,217,2,6,268,0,2,268,1,3,269,1,3,269,2,8,274,2,3,
/* out0010_em-eta10-phi0*/	9,48,1,11,49,2,3,58,0,1,216,0,9,216,1,8,217,0,8,217,2,5,268,0,12,268,1,1,
/* out0011_em-eta11-phi0*/	11,19,5,1,48,0,16,48,1,1,48,2,10,216,0,6,216,1,2,216,2,5,267,0,2,267,1,1,268,0,2,268,2,2,
/* out0012_em-eta12-phi0*/	12,6,3,10,7,2,16,7,3,16,7,4,2,18,5,2,19,5,2,48,2,2,215,0,8,215,1,6,216,0,1,216,2,4,267,0,9,
/* out0013_em-eta13-phi0*/	11,6,0,1,6,1,3,6,2,15,6,3,5,7,0,2,7,4,14,215,0,6,215,1,2,215,2,1,267,0,3,267,2,1,
/* out0014_em-eta14-phi0*/	9,6,1,8,6,2,1,7,0,14,7,1,12,214,0,1,214,1,1,215,0,2,215,2,5,266,0,5,
/* out0015_em-eta15-phi0*/	9,2,3,5,3,2,16,3,3,16,3,4,12,6,4,16,7,1,4,214,0,3,214,1,4,266,0,5,
/* out0016_em-eta16-phi0*/	8,2,2,11,2,3,2,3,0,1,3,4,4,214,0,5,214,2,1,265,0,1,266,0,1,
/* out0017_em-eta17-phi0*/	7,2,1,3,2,2,5,3,0,15,3,1,5,214,0,2,214,2,3,265,0,3,
/* out0018_em-eta18-phi0*/	6,0,4,3,1,1,1,2,4,16,3,1,10,214,0,5,265,0,1,
/* out0019_em-eta19-phi0*/	4,0,4,5,0,5,1,1,0,8,1,1,15,
/* out0020_em-eta0-phi1*/	1,277,3,4,
/* out0021_em-eta1-phi1*/	2,277,2,6,277,3,12,
/* out0022_em-eta2-phi1*/	7,63,1,10,63,2,1,75,1,2,76,1,8,76,2,14,276,3,7,277,2,10,
/* out0023_em-eta3-phi1*/	9,62,1,12,62,2,1,63,2,10,74,1,1,75,0,16,75,1,4,75,2,4,276,2,9,276,3,9,
/* out0024_em-eta4-phi1*/	6,61,1,10,62,2,13,74,0,14,74,1,1,275,3,10,276,2,7,
/* out0025_em-eta5-phi1*/	7,60,1,4,61,0,2,61,1,4,61,2,15,73,0,6,275,2,11,275,3,6,
/* out0026_em-eta6-phi1*/	6,60,0,4,60,1,11,60,2,10,73,0,1,274,5,12,275,2,5,
/* out0027_em-eta7-phi1*/	7,59,0,3,59,1,12,60,0,1,60,2,5,72,0,1,274,4,13,274,5,4,
/* out0028_em-eta8-phi1*/	13,49,1,1,58,1,1,59,0,6,59,1,1,59,2,11,213,1,1,213,2,11,217,1,1,263,0,1,269,1,3,269,2,3,274,3,13,274,4,3,
/* out0029_em-eta9-phi1*/	14,49,1,2,49,2,1,58,0,7,58,1,7,212,0,5,212,1,3,213,1,3,213,2,2,217,1,3,217,2,4,263,0,7,268,1,5,269,1,10,274,3,3,
/* out0030_em-eta10-phi1*/	10,19,2,1,48,1,1,48,2,2,58,0,6,58,2,5,212,0,10,216,1,4,217,2,1,268,1,7,268,2,8,
/* out0031_em-eta11-phi1*/	14,19,2,15,19,3,3,19,4,7,19,5,10,48,1,1,48,2,2,211,0,3,211,1,1,212,2,1,216,1,2,216,2,6,261,0,1,267,1,7,268,2,5,
/* out0032_em-eta12-phi1*/	13,6,0,1,6,3,1,18,4,5,18,5,14,19,0,7,19,4,2,19,5,3,211,0,5,215,1,4,216,2,1,267,0,2,267,1,5,267,2,4,
/* out0033_em-eta13-phi1*/	8,6,0,13,6,1,1,17,2,7,18,4,7,215,1,4,215,2,5,266,1,3,267,2,6,
/* out0034_em-eta14-phi1*/	10,6,0,1,6,1,4,16,5,1,17,2,3,17,5,15,210,0,2,214,1,1,215,2,5,266,0,2,266,1,5,
/* out0035_em-eta15-phi1*/	7,2,0,1,2,3,6,16,4,2,16,5,12,214,1,6,266,0,3,266,2,4,
/* out0036_em-eta16-phi1*/	9,2,0,11,2,1,1,2,3,3,16,4,1,214,1,1,214,2,4,265,0,1,265,1,3,266,2,3,
/* out0037_em-eta17-phi1*/	7,2,0,3,2,1,8,5,2,1,5,5,1,214,2,4,265,0,5,265,1,1,
/* out0038_em-eta18-phi1*/	6,0,4,1,2,1,4,3,1,1,4,5,2,5,5,4,265,0,1,
/* out0039_em-eta19-phi1*/	4,0,4,7,0,5,7,1,0,8,4,5,1,
/* out0040_em-eta0-phi2*/	1,281,0,4,
/* out0041_em-eta1-phi2*/	2,281,0,12,281,1,6,
/* out0042_em-eta2-phi2*/	8,75,1,2,76,1,8,76,2,2,115,0,14,115,1,12,115,2,5,280,0,7,281,1,10,
/* out0043_em-eta3-phi2*/	9,74,1,3,75,1,8,75,2,12,114,0,13,114,1,5,115,0,2,115,2,4,280,0,9,280,1,9,
/* out0044_em-eta4-phi2*/	8,74,0,2,74,1,11,74,2,15,113,0,6,114,0,3,114,2,1,279,0,10,280,1,7,
/* out0045_em-eta5-phi2*/	7,73,0,7,73,1,15,73,2,7,74,2,1,113,0,1,279,0,6,279,1,11,
/* out0046_em-eta6-phi2*/	8,60,1,1,60,2,1,72,0,5,72,1,10,73,0,2,73,2,7,278,0,12,279,1,5,
/* out0047_em-eta7-phi2*/	6,59,1,3,71,1,1,72,0,10,72,2,6,278,0,4,278,1,13,
/* out0048_em-eta8-phi2*/	11,58,1,1,59,2,5,71,0,10,71,1,2,207,0,1,207,2,5,213,1,9,213,2,3,263,1,8,278,1,3,278,2,13,
/* out0049_em-eta9-phi2*/	11,58,1,7,58,2,3,70,0,1,71,0,4,207,2,5,212,1,12,213,1,3,263,0,7,263,1,5,263,2,7,278,2,3,
/* out0050_em-eta10-phi2*/	12,18,3,1,19,3,4,58,2,8,70,0,3,212,0,1,212,1,1,212,2,13,261,0,4,261,1,7,263,0,1,263,2,3,268,2,1,
/* out0051_em-eta11-phi2*/	11,18,0,1,18,2,9,18,3,15,19,3,9,19,4,6,211,0,2,211,1,10,212,2,1,261,0,10,261,2,2,267,1,1,
/* out0052_em-eta12-phi2*/	14,18,1,7,18,2,7,18,4,1,19,0,9,19,1,10,19,4,1,211,0,5,211,2,5,260,0,3,260,1,1,261,0,1,261,2,1,267,1,2,267,2,3,
/* out0053_em-eta13-phi2*/	12,17,2,6,17,3,13,17,4,1,18,4,3,19,1,5,210,0,2,210,1,4,211,0,1,211,2,2,260,0,6,266,1,2,267,2,2,
/* out0054_em-eta14-phi2*/	9,16,2,3,17,0,4,17,3,1,17,4,15,17,5,1,210,0,7,260,0,1,266,1,6,266,2,1,
/* out0055_em-eta15-phi2*/	8,16,4,4,16,5,3,17,0,9,17,1,3,210,0,4,210,2,1,214,1,2,266,2,6,
/* out0056_em-eta16-phi2*/	8,2,0,1,5,2,7,16,4,8,209,1,2,214,1,1,214,2,3,265,1,5,266,2,2,
/* out0057_em-eta17-phi2*/	8,5,2,7,5,4,1,5,5,6,209,0,1,209,1,2,214,2,1,265,0,3,265,1,3,
/* out0058_em-eta18-phi2*/	4,4,5,4,5,0,1,5,4,2,5,5,5,
/* out0059_em-eta19-phi2*/	3,0,5,8,4,4,2,4,5,7,
/* out0060_em-eta0-phi3*/	1,281,3,4,
/* out0061_em-eta1-phi3*/	2,281,2,6,281,3,12,
/* out0062_em-eta2-phi3*/	8,115,1,4,115,2,6,126,0,8,126,1,11,126,2,1,128,2,3,280,3,7,281,2,10,
/* out0063_em-eta3-phi3*/	9,114,1,11,114,2,11,115,2,1,124,0,6,124,1,2,126,0,8,126,2,5,280,2,9,280,3,9,
/* out0064_em-eta4-phi3*/	7,113,0,5,113,1,16,113,2,7,114,2,4,124,0,6,279,3,10,280,2,7,
/* out0065_em-eta5-phi3*/	8,73,1,1,73,2,2,112,0,6,112,1,10,113,0,4,113,2,8,279,2,11,279,3,6,
/* out0066_em-eta6-phi3*/	8,72,1,6,72,2,2,111,0,1,111,1,2,112,0,10,112,2,5,278,5,12,279,2,5,
/* out0067_em-eta7-phi3*/	5,71,1,4,72,2,8,111,0,9,278,4,13,278,5,4,
/* out0068_em-eta8-phi3*/	9,71,0,2,71,1,9,71,2,7,207,0,14,207,1,1,207,2,1,263,1,1,278,3,13,278,4,3,
/* out0069_em-eta9-phi3*/	11,70,0,1,70,1,7,71,2,7,206,1,3,207,1,10,207,2,5,263,1,2,263,2,5,264,1,8,264,2,4,278,3,3,
/* out0070_em-eta10-phi3*/	10,70,0,8,70,1,3,70,2,2,206,0,11,206,1,3,212,2,1,261,1,9,261,2,1,263,2,1,264,1,6,
/* out0071_em-eta11-phi3*/	10,18,0,11,21,2,7,70,0,3,70,2,2,206,0,5,206,2,1,211,1,5,211,2,1,261,2,11,262,1,1,
/* out0072_em-eta12-phi3*/	10,18,0,4,18,1,9,20,5,1,21,2,6,21,5,15,205,0,4,211,2,7,260,0,1,260,1,10,261,2,1,
/* out0073_em-eta13-phi3*/	12,16,0,2,16,3,12,17,3,2,19,1,1,20,4,1,20,5,10,205,0,1,210,1,8,211,2,1,260,0,4,260,1,1,260,2,4,
/* out0074_em-eta14-phi3*/	11,16,0,5,16,1,4,16,2,11,16,3,4,210,0,1,210,1,2,210,2,4,259,0,1,259,1,2,260,0,1,260,2,3,
/* out0075_em-eta15-phi3*/	7,16,1,7,16,2,2,17,0,3,17,1,9,209,1,1,210,2,5,259,0,6,
/* out0076_em-eta16-phi3*/	7,5,2,1,5,3,11,16,4,1,17,1,4,209,1,5,259,0,5,265,1,1,
/* out0077_em-eta17-phi3*/	7,4,2,1,5,3,3,5,4,10,209,0,3,209,1,2,265,0,1,265,1,3,
/* out0078_em-eta18-phi3*/	4,4,2,1,5,0,8,5,4,3,209,0,2,
/* out0079_em-eta19-phi3*/	4,4,4,4,4,5,2,5,0,3,5,1,2,
/* out0080_em-eta0-phi4*/	1,285,0,4,
/* out0081_em-eta1-phi4*/	2,285,0,12,285,1,6,
/* out0082_em-eta2-phi4*/	9,126,1,5,126,2,4,127,1,3,127,2,10,128,0,16,128,1,16,128,2,13,284,0,7,285,1,10,
/* out0083_em-eta3-phi4*/	10,124,0,1,124,1,14,124,2,5,125,1,2,125,2,1,126,2,6,127,0,4,127,1,13,284,0,9,284,1,9,
/* out0084_em-eta4-phi4*/	9,113,2,1,123,0,5,123,1,14,123,2,1,124,0,3,124,2,11,125,1,4,283,0,10,284,1,7,
/* out0085_em-eta5-phi4*/	8,112,1,6,112,2,3,122,0,2,122,1,3,123,0,11,123,2,7,283,0,6,283,1,11,
/* out0086_em-eta6-phi4*/	5,111,1,9,112,2,8,122,0,9,282,0,12,283,1,5,
/* out0087_em-eta7-phi4*/	5,111,0,5,111,1,5,111,2,11,282,0,4,282,1,13,
/* out0088_em-eta8-phi4*/	12,71,2,2,110,0,6,110,1,7,111,0,1,111,2,2,207,0,1,207,1,2,208,0,5,208,2,2,264,2,1,282,1,3,282,2,13,
/* out0089_em-eta9-phi4*/	10,70,1,4,110,0,10,206,1,3,207,1,3,208,0,2,208,2,14,264,0,6,264,1,1,264,2,11,282,2,3,
/* out0090_em-eta10-phi4*/	8,70,1,2,70,2,8,163,1,1,206,1,7,206,2,9,262,2,5,264,0,9,264,1,1,
/* out0091_em-eta11-phi4*/	9,20,3,6,21,2,3,21,3,15,21,4,1,70,2,4,205,1,6,206,2,6,262,1,10,262,2,3,
/* out0092_em-eta12-phi4*/	12,20,2,8,21,0,8,21,3,1,21,4,15,21,5,1,205,0,7,205,1,3,205,2,1,260,1,4,260,2,1,262,0,1,262,1,5,
/* out0093_em-eta13-phi4*/	9,20,4,13,20,5,5,21,0,6,21,1,3,205,0,4,205,2,2,210,1,2,260,2,7,270,1,2,
/* out0094_em-eta14-phi4*/	9,16,0,9,20,4,1,28,5,8,29,5,3,199,1,3,210,2,4,259,1,6,260,2,1,270,1,1,
/* out0095_em-eta15-phi4*/	10,16,1,5,28,4,9,28,5,3,199,1,2,209,1,1,209,2,1,210,2,2,259,0,1,259,1,4,259,2,1,
/* out0096_em-eta16-phi4*/	7,4,3,10,5,3,2,28,4,4,209,1,2,209,2,3,259,0,2,259,2,4,
/* out0097_em-eta17-phi4*/	7,4,2,7,4,3,6,209,0,5,209,1,1,209,2,1,259,0,1,259,2,1,
/* out0098_em-eta18-phi4*/	4,4,1,2,4,2,7,5,0,3,209,0,3,
/* out0099_em-eta19-phi4*/	3,4,4,10,5,0,1,5,1,9,
/* out0100_em-eta0-phi5*/	1,285,3,4,
/* out0101_em-eta1-phi5*/	2,285,2,6,285,3,12,
/* out0102_em-eta2-phi5*/	6,127,0,2,127,2,6,138,0,6,138,2,1,284,3,7,285,2,10,
/* out0103_em-eta3-phi5*/	9,125,0,3,125,1,2,125,2,15,127,0,10,138,0,3,138,1,1,138,2,15,284,2,9,284,3,9,
/* out0104_em-eta4-phi5*/	8,123,1,2,123,2,3,125,0,13,125,1,8,136,1,3,136,2,8,283,3,10,284,2,7,
/* out0105_em-eta5-phi5*/	6,122,1,12,122,2,1,123,2,5,136,1,13,283,2,11,283,3,6,
/* out0106_em-eta6-phi5*/	6,122,0,5,122,1,1,122,2,15,146,2,3,282,5,12,283,2,5,
/* out0107_em-eta7-phi5*/	5,111,2,3,146,1,13,146,2,4,282,4,13,282,5,4,
/* out0108_em-eta8-phi5*/	7,110,1,9,110,2,5,146,1,3,208,0,7,208,1,1,282,3,13,282,4,3,
/* out0109_em-eta9-phi5*/	9,110,2,11,163,2,3,201,1,1,208,0,2,208,1,14,264,0,1,272,0,6,272,1,8,282,3,3,
/* out0110_em-eta10-phi5*/	7,163,1,8,163,2,4,201,0,7,201,1,7,208,1,1,262,2,5,272,0,10,
/* out0111_em-eta11-phi5*/	7,20,0,5,20,3,8,163,1,7,201,0,9,205,1,4,262,0,10,262,2,3,
/* out0112_em-eta12-phi5*/	9,20,0,11,20,1,11,20,2,8,20,3,2,21,0,1,205,1,3,205,2,8,262,0,5,270,2,6,
/* out0113_em-eta13-phi5*/	10,20,1,5,20,4,1,21,0,1,21,1,13,29,2,6,29,5,1,199,2,4,205,2,5,270,1,8,270,2,2,
/* out0114_em-eta14-phi5*/	9,28,5,2,29,0,2,29,2,1,29,4,7,29,5,12,199,1,4,199,2,4,259,1,2,270,1,5,
/* out0115_em-eta15-phi5*/	7,28,4,1,28,5,3,29,0,13,29,1,2,199,1,6,259,1,2,259,2,5,
/* out0116_em-eta16-phi5*/	6,4,0,2,28,4,2,29,1,13,199,1,1,209,2,5,259,2,5,
/* out0117_em-eta17-phi5*/	3,4,0,12,4,1,1,209,2,5,
/* out0118_em-eta18-phi5*/	4,4,0,2,4,1,9,209,0,2,209,2,1,
/* out0119_em-eta19-phi5*/	2,4,1,4,5,1,5,
/* out0120_em-eta0-phi6*/	1,289,0,4,
/* out0121_em-eta1-phi6*/	2,289,0,12,289,1,6,
/* out0122_em-eta2-phi6*/	6,138,0,6,138,1,1,139,1,2,139,2,6,288,0,7,289,1,10,
/* out0123_em-eta3-phi6*/	8,137,0,2,137,1,3,137,2,15,138,0,1,138,1,14,139,1,10,288,0,9,288,1,9,
/* out0124_em-eta4-phi6*/	8,136,0,3,136,2,8,137,0,8,137,1,13,148,1,3,148,2,2,287,0,10,288,1,7,
/* out0125_em-eta5-phi6*/	6,136,0,13,147,1,1,147,2,12,148,1,5,287,0,6,287,1,11,
/* out0126_em-eta6-phi6*/	6,146,2,4,147,0,5,147,1,15,147,2,1,286,0,12,287,1,5,
/* out0127_em-eta7-phi6*/	5,146,0,13,146,2,5,165,1,3,286,0,4,286,1,13,
/* out0128_em-eta8-phi6*/	7,146,0,3,164,1,5,164,2,9,203,0,8,203,2,1,286,1,3,286,2,13,
/* out0129_em-eta9-phi6*/	10,163,2,4,164,1,11,201,1,1,203,0,4,203,1,3,203,2,14,272,1,8,272,2,5,273,1,1,286,2,3,
/* out0130_em-eta10-phi6*/	7,163,0,7,163,2,5,201,1,7,201,2,7,203,2,1,271,2,5,272,2,11,
/* out0131_em-eta11-phi6*/	7,31,2,3,31,5,9,163,0,7,200,2,4,201,2,9,271,1,10,271,2,3,
/* out0132_em-eta12-phi6*/	9,30,4,3,30,5,16,31,0,6,31,4,2,31,5,6,200,1,8,200,2,3,270,2,6,271,1,5,
/* out0133_em-eta13-phi6*/	9,29,2,7,29,3,1,30,4,13,31,0,1,31,1,6,199,2,4,200,1,5,270,0,7,270,2,2,
/* out0134_em-eta14-phi6*/	9,28,2,2,28,3,1,29,2,2,29,3,11,29,4,8,199,0,4,199,2,4,255,2,2,270,0,5,
/* out0135_em-eta15-phi6*/	9,28,0,1,28,1,2,28,2,14,28,3,2,29,0,1,29,4,1,199,0,6,255,1,5,255,2,2,
/* out0136_em-eta16-phi6*/	6,28,1,13,29,1,1,37,5,2,194,1,4,199,0,1,255,1,5,
/* out0137_em-eta17-phi6*/	4,28,1,1,36,5,7,37,5,6,194,1,4,
/* out0138_em-eta18-phi6*/	4,36,4,4,36,5,7,194,0,2,194,1,1,
/* out0139_em-eta19-phi6*/	1,36,4,9,
/* out0140_em-eta0-phi7*/	1,289,3,4,
/* out0141_em-eta1-phi7*/	2,289,2,6,289,3,12,
/* out0142_em-eta2-phi7*/	9,139,0,3,139,2,10,140,0,16,140,1,16,140,2,15,150,1,4,150,2,5,288,3,7,289,2,10,
/* out0143_em-eta3-phi7*/	10,137,0,2,137,2,1,139,0,13,139,1,4,149,0,2,149,1,5,149,2,14,150,1,6,288,2,9,288,3,9,
/* out0144_em-eta4-phi7*/	9,137,0,4,148,0,5,148,1,1,148,2,14,149,0,3,149,1,11,167,1,1,287,3,10,288,2,7,
/* out0145_em-eta5-phi7*/	8,147,0,2,147,2,3,148,0,11,148,1,7,166,1,3,166,2,6,287,2,11,287,3,6,
/* out0146_em-eta6-phi7*/	5,147,0,9,165,2,9,166,1,8,286,5,12,287,2,5,
/* out0147_em-eta7-phi7*/	5,165,0,5,165,1,11,165,2,5,286,4,13,286,5,4,
/* out0148_em-eta8-phi7*/	12,85,1,2,164,0,6,164,2,7,165,0,1,165,1,2,203,0,4,203,1,2,204,0,1,204,2,2,273,2,1,286,3,13,286,4,3,
/* out0149_em-eta9-phi7*/	9,84,2,5,164,0,10,202,2,3,203,1,11,204,2,3,273,0,1,273,1,6,273,2,11,286,3,3,
/* out0150_em-eta10-phi7*/	9,84,1,9,84,2,2,163,0,1,202,1,9,202,2,7,271,0,1,271,2,5,273,0,1,273,1,9,
/* out0151_em-eta11-phi7*/	10,31,2,13,31,3,10,31,4,1,31,5,1,84,1,3,163,0,1,200,2,6,202,1,6,271,0,10,271,2,3,
/* out0152_em-eta12-phi7*/	12,30,2,13,30,3,1,31,0,6,31,3,2,31,4,13,200,0,7,200,1,1,200,2,3,256,1,1,256,2,4,271,0,4,271,1,1,
/* out0153_em-eta13-phi7*/	9,30,1,12,30,2,3,31,0,3,31,1,9,195,2,2,200,0,4,200,1,2,256,1,7,270,0,3,
/* out0154_em-eta14-phi7*/	11,28,3,9,29,3,4,30,1,1,31,1,1,38,5,7,39,5,3,195,1,4,199,0,3,255,2,6,256,1,1,270,0,1,
/* out0155_em-eta15-phi7*/	11,28,0,10,28,3,4,38,4,4,38,5,1,194,1,1,194,2,1,195,1,2,199,0,2,255,0,1,255,1,1,255,2,4,
/* out0156_em-eta16-phi7*/	7,28,0,5,37,2,10,37,5,2,194,1,4,194,2,1,255,0,2,255,1,4,
/* out0157_em-eta17-phi7*/	7,37,0,1,37,4,6,37,5,6,194,0,3,194,1,2,255,0,1,255,1,1,
/* out0158_em-eta18-phi7*/	4,36,5,2,37,0,9,37,1,7,194,0,3,
/* out0159_em-eta19-phi7*/	3,36,4,3,37,0,1,37,1,6,
/* out0160_em-eta0-phi8*/	1,293,0,4,
/* out0161_em-eta1-phi8*/	2,293,0,12,293,1,6,
/* out0162_em-eta2-phi8*/	8,140,2,1,150,0,8,150,1,1,150,2,11,169,1,6,169,2,4,292,0,7,293,1,10,
/* out0163_em-eta3-phi8*/	9,149,0,6,149,2,2,150,0,8,150,1,5,168,1,11,168,2,11,169,1,1,292,0,9,292,1,9,
/* out0164_em-eta4-phi8*/	7,149,0,5,167,0,5,167,1,7,167,2,16,168,1,4,291,0,10,292,1,7,
/* out0165_em-eta5-phi8*/	8,87,1,2,87,2,1,166,0,6,166,2,10,167,0,4,167,1,8,291,0,6,291,1,11,
/* out0166_em-eta6-phi8*/	8,86,1,2,86,2,6,165,0,1,165,2,2,166,0,10,166,1,5,290,0,12,291,1,5,
/* out0167_em-eta7-phi8*/	5,85,2,4,86,1,8,165,0,9,290,0,4,290,1,13,
/* out0168_em-eta8-phi8*/	9,85,0,2,85,1,7,85,2,9,204,0,14,204,1,2,204,2,1,258,2,1,290,1,3,290,2,13,
/* out0169_em-eta9-phi8*/	11,84,0,1,84,2,7,85,1,7,202,2,3,204,1,6,204,2,10,258,1,5,258,2,2,273,0,8,273,2,4,290,2,3,
/* out0170_em-eta10-phi8*/	10,84,0,8,84,1,2,84,2,2,197,1,1,202,0,11,202,2,3,257,1,1,257,2,9,258,1,1,273,0,6,
/* out0171_em-eta11-phi8*/	12,30,3,2,31,3,4,40,5,4,41,5,7,84,0,3,84,1,2,196,1,1,196,2,5,202,0,5,202,1,1,257,1,11,271,0,1,
/* out0172_em-eta12-phi8*/	9,30,0,8,30,3,13,40,4,5,40,5,7,196,1,7,200,0,4,256,0,1,256,2,10,257,1,1,
/* out0173_em-eta13-phi8*/	11,30,0,8,30,1,3,39,2,10,39,5,6,40,4,1,195,2,8,196,1,1,200,0,1,256,0,4,256,1,4,256,2,1,
/* out0174_em-eta14-phi8*/	11,38,5,5,39,0,5,39,4,6,39,5,7,195,0,1,195,1,4,195,2,2,255,0,1,255,2,2,256,0,1,256,1,3,
/* out0175_em-eta15-phi8*/	7,38,4,9,38,5,3,39,0,4,39,1,4,194,2,1,195,1,5,255,0,6,
/* out0176_em-eta16-phi8*/	7,37,2,6,37,3,6,38,4,3,39,1,2,194,2,6,250,1,1,255,0,5,
/* out0177_em-eta17-phi8*/	6,36,2,2,37,3,3,37,4,9,194,0,5,194,2,2,250,1,4,
/* out0178_em-eta18-phi8*/	5,36,1,3,36,2,8,37,0,3,37,4,1,194,0,2,
/* out0179_em-eta19-phi8*/	4,36,1,4,36,2,2,37,0,2,37,1,3,
/* out0180_em-eta0-phi9*/	1,293,3,4,
/* out0181_em-eta1-phi9*/	2,293,2,6,293,3,12,
/* out0182_em-eta2-phi9*/	8,89,2,2,90,0,2,90,1,8,169,0,14,169,1,5,169,2,12,292,3,7,293,2,10,
/* out0183_em-eta3-phi9*/	9,88,2,3,89,1,12,89,2,8,168,0,13,168,2,5,169,0,2,169,1,4,292,2,9,292,3,9,
/* out0184_em-eta4-phi9*/	8,88,0,2,88,1,15,88,2,11,167,0,6,168,0,3,168,1,1,291,3,10,292,2,7,
/* out0185_em-eta5-phi9*/	7,87,0,7,87,1,7,87,2,15,88,1,1,167,0,1,291,2,11,291,3,6,
/* out0186_em-eta6-phi9*/	8,86,0,5,86,2,10,87,0,2,87,1,7,100,1,1,100,2,1,290,5,12,291,2,5,
/* out0187_em-eta7-phi9*/	6,85,2,1,86,0,10,86,1,6,99,2,3,290,4,13,290,5,4,
/* out0188_em-eta8-phi9*/	11,85,0,10,85,2,2,98,2,1,99,1,5,198,0,3,198,1,9,204,0,1,204,1,4,258,2,8,290,3,13,290,4,3,
/* out0189_em-eta9-phi9*/	11,84,0,1,85,0,4,98,1,3,98,2,7,197,2,12,198,1,3,204,1,4,258,0,7,258,1,7,258,2,5,290,3,3,
/* out0190_em-eta10-phi9*/	11,41,2,5,84,0,3,98,1,8,197,0,1,197,1,13,197,2,1,253,1,1,257,0,4,257,2,7,258,0,1,258,1,3,
/* out0191_em-eta11-phi9*/	12,40,5,1,41,0,1,41,2,11,41,3,5,41,4,14,41,5,9,196,0,2,196,2,10,197,1,1,252,2,1,257,0,10,257,1,2,
/* out0192_em-eta12-phi9*/	13,40,2,2,40,4,6,40,5,4,41,0,15,41,1,7,196,0,5,196,1,5,252,1,3,252,2,2,256,0,3,256,2,1,257,0,1,257,1,1,
/* out0193_em-eta13-phi9*/	12,39,2,6,39,3,13,39,4,1,40,4,4,41,1,5,195,0,2,195,2,4,196,0,1,196,1,2,251,2,2,252,1,2,256,0,6,
/* out0194_em-eta14-phi9*/	9,38,2,11,38,3,1,39,0,2,39,3,1,39,4,9,195,0,7,251,1,1,251,2,6,256,0,1,
/* out0195_em-eta15-phi9*/	8,38,1,6,38,2,5,39,0,5,39,1,4,190,2,2,195,0,4,195,1,1,251,1,6,
/* out0196_em-eta16-phi9*/	10,36,3,2,37,3,5,38,1,3,39,1,6,190,1,3,190,2,1,194,2,2,250,1,2,250,2,2,251,1,2,
/* out0197_em-eta17-phi9*/	8,36,2,1,36,3,11,37,3,2,190,1,1,194,0,1,194,2,3,250,1,5,250,2,1,
/* out0198_em-eta18-phi9*/	5,36,0,5,36,1,2,36,2,3,36,3,2,250,1,1,
/* out0199_em-eta19-phi9*/	3,8,3,1,36,0,2,36,1,7,
/* out0200_em-eta0-phi10*/	1,297,0,4,
/* out0201_em-eta1-phi10*/	2,297,0,12,297,1,6,
/* out0202_em-eta2-phi10*/	7,89,2,2,90,0,14,90,1,8,103,1,1,103,2,10,296,0,7,297,1,10,
/* out0203_em-eta3-phi10*/	9,88,2,1,89,0,16,89,1,4,89,2,4,102,1,1,102,2,12,103,1,10,296,0,9,296,1,9,
/* out0204_em-eta4-phi10*/	6,88,0,14,88,2,1,101,2,10,102,1,13,295,0,10,296,1,7,
/* out0205_em-eta5-phi10*/	7,87,0,6,100,2,4,101,0,2,101,1,15,101,2,4,295,0,6,295,1,11,
/* out0206_em-eta6-phi10*/	6,87,0,1,100,0,4,100,1,10,100,2,11,294,0,12,295,1,5,
/* out0207_em-eta7-phi10*/	7,86,0,1,99,0,3,99,2,12,100,0,1,100,1,5,294,0,4,294,1,13,
/* out0208_em-eta8-phi10*/	12,98,2,1,99,0,6,99,1,11,99,2,1,193,2,1,198,0,11,198,1,1,254,0,3,254,1,3,258,0,1,294,1,3,294,2,13,
/* out0209_em-eta9-phi10*/	12,98,0,7,98,2,7,193,1,4,193,2,3,197,0,5,197,2,3,198,0,2,198,1,3,253,2,5,254,1,10,258,0,7,294,2,3,
/* out0210_em-eta10-phi10*/	9,41,3,1,53,0,1,98,0,6,98,1,5,192,2,4,193,1,1,197,0,10,253,1,8,253,2,7,
/* out0211_em-eta11-phi10*/	14,40,0,3,40,2,5,40,3,15,41,3,10,41,4,2,53,0,1,192,1,6,192,2,2,196,0,3,196,2,1,197,1,1,252,2,7,253,1,5,257,0,1,
/* out0212_em-eta12-phi10*/	12,15,5,1,40,0,9,40,1,12,40,2,9,40,3,1,41,1,1,191,2,4,192,1,1,196,0,5,252,0,2,252,1,4,252,2,5,
/* out0213_em-eta13-phi10*/	10,14,5,7,15,5,6,38,3,5,39,3,2,40,1,4,41,1,3,191,1,5,191,2,4,251,2,3,252,1,6,
/* out0214_em-eta14-phi10*/	9,14,4,2,14,5,2,38,0,9,38,3,10,190,2,1,191,1,5,195,0,2,251,0,2,251,2,5,
/* out0215_em-eta15-phi10*/	7,13,2,3,13,5,2,38,0,7,38,1,6,190,2,6,251,0,3,251,1,4,
/* out0216_em-eta16-phi10*/	7,12,5,5,13,5,10,38,1,1,190,1,4,190,2,1,250,2,4,251,1,3,
/* out0217_em-eta17-phi10*/	7,12,4,3,12,5,8,36,0,1,36,3,1,190,1,4,250,1,1,250,2,5,
/* out0218_em-eta18-phi10*/	4,8,0,1,12,4,4,36,0,6,250,1,1,
/* out0219_em-eta19-phi10*/	3,8,0,6,8,3,13,36,0,2,
/* out0220_em-eta0-phi11*/	1,297,3,4,
/* out0221_em-eta1-phi11*/	2,297,2,6,297,3,12,
/* out0222_em-eta2-phi11*/	4,103,0,8,103,2,6,296,3,7,297,2,10,
/* out0223_em-eta3-phi11*/	6,102,0,7,102,2,4,103,0,8,103,1,5,296,2,9,296,3,9,
/* out0224_em-eta4-phi11*/	9,57,0,15,57,1,4,57,2,1,101,0,3,101,2,2,102,0,9,102,1,2,295,3,10,296,2,7,
/* out0225_em-eta5-phi11*/	8,56,0,10,56,1,4,57,0,1,57,2,3,101,0,11,101,1,1,295,2,11,295,3,6,
/* out0226_em-eta6-phi11*/	7,55,0,3,55,1,3,56,0,6,56,2,4,100,0,10,294,5,12,295,2,5,
/* out0227_em-eta7-phi11*/	7,55,0,13,55,1,1,55,2,2,99,0,3,100,0,1,294,4,13,294,5,4,
/* out0228_em-eta8-phi11*/	9,54,0,7,54,1,4,55,2,1,99,0,4,193,0,1,193,2,7,254,0,5,294,3,13,294,4,3,
/* out0229_em-eta9-phi11*/	12,54,0,9,54,2,4,98,0,2,193,0,7,193,1,6,193,2,5,249,0,6,253,0,2,253,2,3,254,0,8,254,1,3,294,3,3,
/* out0230_em-eta10-phi11*/	11,53,0,7,53,1,4,98,0,1,192,0,2,192,2,8,193,0,1,193,1,5,248,0,1,249,0,1,253,0,12,253,2,1,
/* out0231_em-eta11-phi11*/	11,40,0,1,53,0,7,53,2,2,192,0,6,192,1,5,192,2,2,248,0,6,252,0,2,252,2,1,253,0,2,253,1,2,
/* out0232_em-eta12-phi11*/	12,15,2,16,15,3,4,15,4,2,15,5,3,40,0,3,53,2,2,191,0,1,191,2,6,192,0,1,192,1,4,248,0,1,252,0,9,
/* out0233_em-eta13-phi11*/	10,14,5,4,15,0,8,15,4,10,15,5,6,191,0,5,191,1,1,191,2,2,247,0,5,252,0,3,252,1,1,
/* out0234_em-eta14-phi11*/	9,14,4,13,14,5,3,15,0,3,15,1,4,190,2,1,191,0,2,191,1,5,247,0,2,251,0,5,
/* out0235_em-eta15-phi11*/	9,13,2,13,13,3,4,13,4,1,13,5,1,14,4,1,190,0,3,190,2,4,246,0,2,251,0,5,
/* out0236_em-eta16-phi11*/	7,13,0,4,13,4,11,13,5,3,190,0,4,190,1,1,246,0,4,251,0,1,
/* out0237_em-eta17-phi11*/	8,12,4,2,12,5,3,13,0,8,13,1,2,190,0,2,190,1,3,246,0,2,250,2,3,
/* out0238_em-eta18-phi11*/	5,8,0,3,12,4,7,13,1,2,250,1,1,250,2,1,
/* out0239_em-eta19-phi11*/	4,8,0,6,8,1,3,8,2,11,8,3,2,
/* out0240_em-eta0-phi12*/	1,301,0,4,
/* out0241_em-eta1-phi12*/	2,301,0,12,301,1,6,
/* out0242_em-eta2-phi12*/	4,69,0,8,69,1,6,300,0,7,301,1,10,
/* out0243_em-eta3-phi12*/	6,68,0,7,68,1,4,69,0,8,69,2,5,300,0,9,300,1,9,
/* out0244_em-eta4-phi12*/	8,57,1,12,57,2,8,67,0,3,67,1,2,68,0,9,68,2,2,299,0,10,300,1,7,
/* out0245_em-eta5-phi12*/	7,56,1,12,56,2,2,57,2,4,67,0,11,67,2,1,299,0,6,299,1,11,
/* out0246_em-eta6-phi12*/	5,55,1,6,56,2,10,66,0,10,298,0,12,299,1,5,
/* out0247_em-eta7-phi12*/	6,55,1,6,55,2,11,65,0,3,66,0,1,298,0,4,298,1,13,
/* out0248_em-eta8-phi12*/	8,54,1,11,55,2,2,65,0,4,189,0,9,193,0,1,249,1,3,298,1,3,298,2,13,
/* out0249_em-eta9-phi12*/	12,54,1,1,54,2,12,64,0,2,188,0,3,188,1,3,189,0,4,189,2,3,193,0,6,249,0,7,249,1,9,249,2,4,298,2,3,
/* out0250_em-eta10-phi12*/	9,53,1,11,64,0,1,188,0,12,188,2,1,192,0,2,248,0,1,248,1,6,249,0,2,249,2,7,
/* out0251_em-eta11-phi12*/	10,27,5,1,53,2,9,187,0,4,187,1,2,188,0,1,188,2,1,192,0,5,248,0,6,248,1,4,248,2,3,
/* out0252_em-eta12-phi12*/	12,14,3,10,15,3,12,15,4,1,26,5,2,27,5,2,53,2,2,187,0,9,191,0,1,247,0,1,247,1,4,248,0,1,248,2,5,
/* out0253_em-eta13-phi12*/	13,14,0,1,14,1,3,14,2,15,14,3,5,15,0,2,15,4,3,186,0,1,187,0,1,187,2,1,191,0,5,247,0,5,247,1,3,247,2,1,
/* out0254_em-eta14-phi12*/	8,14,1,8,14,2,1,15,0,3,15,1,11,186,0,6,191,0,2,247,0,3,247,2,5,
/* out0255_em-eta15-phi12*/	9,12,3,5,13,3,12,13,4,1,15,1,1,186,0,4,190,0,2,246,0,2,246,1,4,247,2,1,
/* out0256_em-eta16-phi12*/	7,12,2,11,12,3,2,13,4,3,185,0,1,190,0,4,246,0,4,246,1,1,
/* out0257_em-eta17-phi12*/	8,12,1,3,12,2,5,13,0,4,13,1,2,185,0,3,190,0,1,246,0,2,246,2,2,
/* out0258_em-eta18-phi12*/	4,8,1,4,13,1,9,185,1,1,246,2,1,
/* out0259_em-eta19-phi12*/	5,8,1,8,8,2,5,8,4,12,9,0,16,9,1,5,
/* out0260_em-eta0-phi13*/	1,301,3,4,
/* out0261_em-eta1-phi13*/	2,301,2,6,301,3,12,
/* out0262_em-eta2-phi13*/	7,69,1,10,69,2,1,82,1,2,83,0,14,83,2,8,300,3,7,301,2,10,
/* out0263_em-eta3-phi13*/	9,68,1,12,68,2,1,69,2,10,81,1,1,82,0,16,82,1,4,82,2,4,300,2,9,300,3,9,
/* out0264_em-eta4-phi13*/	6,67,1,10,68,2,13,81,0,14,81,1,1,299,3,10,300,2,7,
/* out0265_em-eta5-phi13*/	7,66,1,4,67,0,2,67,1,4,67,2,15,80,0,6,299,2,11,299,3,6,
/* out0266_em-eta6-phi13*/	6,66,0,4,66,1,11,66,2,10,80,0,1,298,5,12,299,2,5,
/* out0267_em-eta7-phi13*/	7,65,0,3,65,1,12,66,0,1,66,2,5,79,0,1,298,4,13,298,5,4,
/* out0268_em-eta8-phi13*/	10,64,1,1,65,0,6,65,1,1,65,2,11,184,0,2,189,0,3,189,2,7,245,0,7,298,3,13,298,4,3,
/* out0269_em-eta9-phi13*/	12,64,0,7,64,1,7,184,0,6,188,1,9,189,2,6,244,0,2,244,1,3,245,0,6,245,2,4,249,1,4,249,2,3,298,3,3,
/* out0270_em-eta10-phi13*/	9,27,2,1,53,1,1,64,0,6,64,2,5,188,1,4,188,2,11,244,0,12,248,1,2,249,2,2,
/* out0271_em-eta11-phi13*/	13,27,2,15,27,3,3,27,4,7,27,5,10,53,2,1,182,0,1,187,1,9,188,2,2,243,0,2,244,0,1,244,2,1,248,1,4,248,2,5,
/* out0272_em-eta12-phi13*/	13,14,0,1,14,3,1,26,4,5,26,5,14,27,0,7,27,4,2,27,5,3,187,0,2,187,1,2,187,2,6,243,0,6,247,1,3,248,2,3,
/* out0273_em-eta13-phi13*/	9,14,0,13,14,1,1,23,2,7,26,4,7,186,1,5,187,2,4,243,0,1,247,1,6,247,2,3,
/* out0274_em-eta14-phi13*/	10,14,0,1,14,1,4,22,5,1,23,2,3,23,5,15,186,0,3,186,1,4,186,2,1,242,0,1,247,2,6,
/* out0275_em-eta15-phi13*/	8,12,0,1,12,3,6,22,4,2,22,5,12,186,0,2,186,2,4,242,0,1,246,1,6,
/* out0276_em-eta16-phi13*/	8,12,0,11,12,1,1,12,3,3,22,4,1,185,0,5,186,2,1,246,1,3,246,2,3,
/* out0277_em-eta17-phi13*/	7,11,2,1,11,5,1,12,0,3,12,1,8,185,0,4,185,1,2,246,2,5,
/* out0278_em-eta18-phi13*/	7,8,1,1,9,1,1,10,5,2,11,5,4,12,1,4,13,1,1,246,2,1,
/* out0279_em-eta19-phi13*/	3,8,4,3,9,1,10,10,5,1,
/* out0280_em-eta0-phi14*/	1,305,0,4,
/* out0281_em-eta1-phi14*/	2,305,0,12,305,1,6,
/* out0282_em-eta2-phi14*/	8,82,1,2,83,0,2,83,2,8,121,0,14,121,1,12,121,2,5,304,0,7,305,1,10,
/* out0283_em-eta3-phi14*/	9,81,1,3,82,1,8,82,2,12,120,0,13,120,1,5,121,0,2,121,2,4,304,0,9,304,1,9,
/* out0284_em-eta4-phi14*/	8,81,0,2,81,1,11,81,2,15,119,0,6,120,0,3,120,2,1,303,0,10,304,1,7,
/* out0285_em-eta5-phi14*/	7,80,0,7,80,1,15,80,2,7,81,2,1,119,0,1,303,0,6,303,1,11,
/* out0286_em-eta6-phi14*/	8,66,1,1,66,2,1,79,0,5,79,1,10,80,0,2,80,2,7,302,0,12,303,1,5,
/* out0287_em-eta7-phi14*/	6,65,1,3,78,1,1,79,0,10,79,2,6,302,0,4,302,1,13,
/* out0288_em-eta8-phi14*/	12,64,1,1,65,2,5,78,0,10,78,1,2,184,0,1,184,1,12,240,0,1,240,2,3,245,0,3,245,2,5,302,1,3,302,2,13,
/* out0289_em-eta9-phi14*/	11,64,1,7,64,2,3,77,0,1,78,0,4,184,0,7,184,1,2,184,2,10,240,2,7,244,1,8,245,2,7,302,2,3,
/* out0290_em-eta10-phi14*/	11,26,3,1,27,3,4,64,2,8,77,0,3,182,0,7,182,1,7,184,2,1,188,2,1,244,0,1,244,1,4,244,2,11,
/* out0291_em-eta11-phi14*/	11,26,0,1,26,2,9,26,3,15,27,3,9,27,4,6,182,0,8,182,2,3,187,1,2,243,0,1,243,1,9,244,2,3,
/* out0292_em-eta12-phi14*/	13,26,1,7,26,2,7,26,4,1,27,0,9,27,1,10,27,4,1,180,0,4,180,1,1,187,1,1,187,2,4,243,0,5,243,1,2,243,2,4,
/* out0293_em-eta13-phi14*/	12,23,2,6,23,3,13,23,4,1,26,4,3,27,1,5,180,0,6,186,1,3,187,2,1,242,0,1,242,1,3,243,0,1,243,2,3,
/* out0294_em-eta14-phi14*/	9,22,2,3,23,0,4,23,3,1,23,4,15,23,5,1,186,1,4,186,2,3,242,0,7,242,1,1,
/* out0295_em-eta15-phi14*/	7,22,4,4,22,5,3,23,0,9,23,1,3,186,2,6,242,0,5,246,1,1,
/* out0296_em-eta16-phi14*/	9,11,2,7,12,0,1,22,4,8,185,0,3,185,1,3,186,2,1,241,1,1,246,1,1,246,2,2,
/* out0297_em-eta17-phi14*/	6,11,2,7,11,4,1,11,5,6,185,1,5,241,1,3,246,2,2,
/* out0298_em-eta18-phi14*/	5,10,5,4,11,0,1,11,4,2,11,5,5,241,0,1,
/* out0299_em-eta19-phi14*/	3,8,4,1,10,4,2,10,5,7,
/* out0300_em-eta0-phi15*/	1,305,3,4,
/* out0301_em-eta1-phi15*/	2,305,2,6,305,3,12,
/* out0302_em-eta2-phi15*/	8,121,1,4,121,2,6,134,0,8,134,1,11,134,2,1,135,0,1,304,3,7,305,2,10,
/* out0303_em-eta3-phi15*/	9,120,1,11,120,2,11,121,2,1,132,0,6,132,1,2,134,0,8,134,2,5,304,2,9,304,3,9,
/* out0304_em-eta4-phi15*/	7,119,0,5,119,1,16,119,2,7,120,2,4,132,0,6,303,3,10,304,2,7,
/* out0305_em-eta5-phi15*/	8,80,1,1,80,2,2,118,0,6,118,1,10,119,0,4,119,2,8,303,2,11,303,3,6,
/* out0306_em-eta6-phi15*/	8,79,1,6,79,2,2,117,0,1,117,1,2,118,0,10,118,2,5,302,5,12,303,2,5,
/* out0307_em-eta7-phi15*/	5,78,1,4,79,2,8,117,0,9,302,4,13,302,5,4,
/* out0308_em-eta8-phi15*/	8,78,0,2,78,1,9,78,2,7,183,2,2,184,1,2,240,0,11,302,3,13,302,4,3,
/* out0309_em-eta9-phi15*/	10,77,0,1,77,1,7,78,2,7,183,1,10,183,2,2,184,2,5,240,0,3,240,1,11,240,2,6,302,3,3,
/* out0310_em-eta10-phi15*/	10,77,0,8,77,1,3,77,2,2,182,1,9,182,2,3,183,1,3,238,0,8,238,1,6,244,1,1,244,2,1,
/* out0311_em-eta11-phi15*/	10,25,2,7,26,0,11,77,0,3,77,2,2,180,1,2,181,1,1,182,2,10,238,0,8,238,2,1,243,1,4,
/* out0312_em-eta12-phi15*/	10,24,5,1,25,2,6,25,5,15,26,0,4,26,1,9,180,0,1,180,1,9,237,0,3,243,1,1,243,2,7,
/* out0313_em-eta13-phi15*/	11,22,0,2,22,3,12,23,3,2,24,4,1,24,5,10,27,1,1,180,0,4,180,2,5,237,0,2,242,1,6,243,2,2,
/* out0314_em-eta14-phi15*/	11,22,0,5,22,1,4,22,2,11,22,3,4,179,0,2,179,1,3,180,0,1,180,2,2,242,0,1,242,1,4,242,2,3,
/* out0315_em-eta15-phi15*/	6,22,1,7,22,2,2,23,0,3,23,1,9,179,0,6,242,2,6,
/* out0316_em-eta16-phi15*/	7,11,2,1,11,3,11,22,4,1,23,1,4,179,0,4,185,1,2,241,1,5,
/* out0317_em-eta17-phi15*/	6,10,2,1,11,3,3,11,4,10,185,1,3,241,0,2,241,1,3,
/* out0318_em-eta18-phi15*/	4,10,2,1,11,0,8,11,4,3,241,0,3,
/* out0319_em-eta19-phi15*/	4,10,4,4,10,5,2,11,0,3,11,1,2,
/* out0320_em-eta0-phi16*/	1,309,0,4,
/* out0321_em-eta1-phi16*/	2,309,0,12,309,1,6,
/* out0322_em-eta2-phi16*/	9,133,1,3,133,2,10,134,1,5,134,2,4,135,0,15,135,1,16,135,2,16,308,0,7,309,1,10,
/* out0323_em-eta3-phi16*/	10,131,1,2,131,2,1,132,0,1,132,1,14,132,2,5,133,0,4,133,1,13,134,2,6,308,0,9,308,1,9,
/* out0324_em-eta4-phi16*/	9,119,2,1,130,0,5,130,1,14,130,2,1,131,1,4,132,0,3,132,2,11,307,0,10,308,1,7,
/* out0325_em-eta5-phi16*/	8,118,1,6,118,2,3,129,0,2,129,1,3,130,0,11,130,2,7,307,0,6,307,1,11,
/* out0326_em-eta6-phi16*/	5,117,1,9,118,2,8,129,0,9,306,0,12,307,1,5,
/* out0327_em-eta7-phi16*/	5,117,0,5,117,1,5,117,2,11,306,0,4,306,1,13,
/* out0328_em-eta8-phi16*/	11,78,2,2,116,0,6,116,1,7,117,0,1,117,2,2,183,2,4,239,0,3,240,0,1,240,1,1,306,1,3,306,2,13,
/* out0329_em-eta9-phi16*/	10,77,1,4,116,0,10,183,0,9,183,1,2,183,2,8,238,1,1,239,0,4,239,2,14,240,1,4,306,2,3,
/* out0330_em-eta10-phi16*/	10,77,1,2,77,2,8,156,1,1,181,1,2,181,2,7,183,0,6,183,1,1,238,1,9,238,2,6,239,2,2,
/* out0331_em-eta11-phi16*/	10,24,3,6,25,2,3,25,3,15,25,4,1,77,2,4,181,0,1,181,1,11,181,2,1,237,1,4,238,2,9,
/* out0332_em-eta12-phi16*/	13,24,2,8,25,0,8,25,3,1,25,4,15,25,5,1,180,1,4,180,2,3,181,0,1,181,1,2,218,1,1,237,0,5,237,1,6,237,2,1,
/* out0333_em-eta13-phi16*/	9,24,4,13,24,5,5,25,0,6,25,1,3,180,2,6,218,1,2,237,0,6,237,2,2,242,1,1,
/* out0334_em-eta14-phi16*/	8,22,0,9,24,4,1,32,5,8,33,5,3,179,1,7,231,1,2,242,1,1,242,2,4,
/* out0335_em-eta15-phi16*/	9,22,1,5,32,4,9,32,5,3,179,0,2,179,1,2,179,2,2,231,1,2,241,1,1,242,2,3,
/* out0336_em-eta16-phi16*/	7,10,3,10,11,3,2,32,4,4,179,0,2,179,2,4,241,1,2,241,2,3,
/* out0337_em-eta17-phi16*/	6,10,2,7,10,3,6,179,2,1,241,0,3,241,1,1,241,2,2,
/* out0338_em-eta18-phi16*/	4,10,1,2,10,2,7,11,0,3,241,0,4,
/* out0339_em-eta19-phi16*/	3,10,4,10,11,0,1,11,1,9,
/* out0340_em-eta0-phi17*/	1,309,3,4,
/* out0341_em-eta1-phi17*/	2,309,2,6,309,3,12,
/* out0342_em-eta2-phi17*/	6,133,0,2,133,2,6,145,0,6,145,2,1,308,3,7,309,2,10,
/* out0343_em-eta3-phi17*/	9,131,0,3,131,1,2,131,2,15,133,0,10,145,0,3,145,1,1,145,2,15,308,2,9,308,3,9,
/* out0344_em-eta4-phi17*/	8,130,1,2,130,2,3,131,0,13,131,1,8,141,1,3,141,2,8,307,3,10,308,2,7,
/* out0345_em-eta5-phi17*/	6,129,1,12,129,2,1,130,2,5,141,1,13,307,2,11,307,3,6,
/* out0346_em-eta6-phi17*/	6,129,0,5,129,1,1,129,2,15,151,2,3,306,5,12,307,2,5,
/* out0347_em-eta7-phi17*/	5,117,2,3,151,1,13,151,2,4,306,4,13,306,5,4,
/* out0348_em-eta8-phi17*/	7,116,1,9,116,2,5,151,1,3,221,1,1,239,0,2,306,3,13,306,4,3,
/* out0349_em-eta9-phi17*/	8,116,2,11,156,2,3,183,0,1,221,0,9,221,1,7,239,0,7,239,1,13,306,3,3,
/* out0350_em-eta10-phi17*/	8,156,1,8,156,2,4,181,0,1,181,2,7,221,0,7,235,0,5,235,1,8,239,1,3,
/* out0351_em-eta11-phi17*/	7,24,0,5,24,3,7,156,1,7,181,0,11,181,2,1,235,0,11,237,1,2,
/* out0352_em-eta12-phi17*/	10,24,0,11,24,1,11,24,2,8,24,3,3,25,0,1,181,0,2,218,1,1,218,2,7,237,1,4,237,2,6,
/* out0353_em-eta13-phi17*/	10,24,1,5,24,4,1,25,0,1,25,1,13,33,2,6,33,5,1,218,1,8,218,2,1,231,2,2,237,2,7,
/* out0354_em-eta14-phi17*/	9,32,5,2,33,0,2,33,2,1,33,4,7,33,5,12,179,1,3,218,1,4,231,1,3,231,2,5,
/* out0355_em-eta15-phi17*/	7,32,4,1,32,5,3,33,0,13,33,1,2,179,1,1,179,2,5,231,1,7,
/* out0356_em-eta16-phi17*/	6,10,0,2,32,4,2,33,1,13,179,2,4,231,1,2,241,2,4,
/* out0357_em-eta17-phi17*/	3,10,0,12,10,1,1,241,2,5,
/* out0358_em-eta18-phi17*/	4,10,0,2,10,1,9,241,0,3,241,2,2,
/* out0359_em-eta19-phi17*/	2,10,1,4,11,1,5,
/* out0360_em-eta0-phi18*/	1,313,0,4,
/* out0361_em-eta1-phi18*/	2,313,0,12,313,1,6,
/* out0362_em-eta2-phi18*/	6,143,1,2,143,2,6,145,0,6,145,1,1,312,0,7,313,1,10,
/* out0363_em-eta3-phi18*/	8,142,0,2,142,1,3,142,2,15,143,1,10,145,0,1,145,1,14,312,0,9,312,1,9,
/* out0364_em-eta4-phi18*/	8,141,0,3,141,2,8,142,0,8,142,1,13,153,1,3,153,2,2,311,0,10,312,1,7,
/* out0365_em-eta5-phi18*/	6,141,0,13,152,1,1,152,2,12,153,1,5,311,0,6,311,1,11,
/* out0366_em-eta6-phi18*/	6,151,2,4,152,0,5,152,1,15,152,2,1,310,0,12,311,1,5,
/* out0367_em-eta7-phi18*/	5,151,0,13,151,2,5,158,1,3,310,0,4,310,1,13,
/* out0368_em-eta8-phi18*/	7,151,0,3,157,1,5,157,2,9,221,1,1,236,0,2,310,1,3,310,2,13,
/* out0369_em-eta9-phi18*/	9,156,2,4,157,1,11,220,1,1,221,1,7,221,2,9,236,0,9,236,1,2,236,2,13,310,2,3,
/* out0370_em-eta10-phi18*/	9,156,0,7,156,2,5,219,1,1,219,2,7,221,2,7,235,1,8,235,2,5,236,1,1,236,2,3,
/* out0371_em-eta11-phi18*/	7,35,2,3,35,5,9,156,0,7,219,1,11,219,2,1,232,2,2,235,2,11,
/* out0372_em-eta12-phi18*/	10,34,4,3,34,5,16,35,0,6,35,4,2,35,5,6,218,0,1,218,2,7,219,1,2,232,1,6,232,2,4,
/* out0373_em-eta13-phi18*/	9,33,2,7,33,3,1,34,4,13,35,0,1,35,1,6,218,0,8,218,2,1,231,2,3,232,1,7,
/* out0374_em-eta14-phi18*/	9,32,2,2,32,3,1,33,2,2,33,3,11,33,4,8,175,2,3,218,0,3,231,0,2,231,2,5,
/* out0375_em-eta15-phi18*/	9,32,0,1,32,1,2,32,2,14,32,3,2,33,0,1,33,4,1,175,1,5,175,2,1,231,0,6,
/* out0376_em-eta16-phi18*/	6,32,1,13,33,1,1,43,5,2,175,1,4,226,1,3,231,0,2,
/* out0377_em-eta17-phi18*/	4,32,1,1,42,5,7,43,5,6,226,1,4,
/* out0378_em-eta18-phi18*/	4,42,4,4,42,5,7,226,0,2,226,1,2,
/* out0379_em-eta19-phi18*/	1,42,4,9,
/* out0380_em-eta0-phi19*/	1,313,3,4,
/* out0381_em-eta1-phi19*/	2,313,2,6,313,3,12,
/* out0382_em-eta2-phi19*/	9,143,0,3,143,2,10,144,0,16,144,1,16,144,2,15,155,1,4,155,2,5,312,3,7,313,2,10,
/* out0383_em-eta3-phi19*/	10,142,0,2,142,2,1,143,0,13,143,1,4,154,0,1,154,1,5,154,2,14,155,1,6,312,2,9,312,3,9,
/* out0384_em-eta4-phi19*/	9,142,0,4,153,0,5,153,1,1,153,2,14,154,0,3,154,1,11,160,1,1,311,3,10,312,2,7,
/* out0385_em-eta5-phi19*/	8,152,0,2,152,2,3,153,0,11,153,1,7,159,1,3,159,2,6,311,2,11,311,3,6,
/* out0386_em-eta6-phi19*/	5,152,0,9,158,2,9,159,1,8,310,5,12,311,2,5,
/* out0387_em-eta7-phi19*/	5,158,0,5,158,1,11,158,2,5,310,4,13,310,5,4,
/* out0388_em-eta8-phi19*/	11,92,1,2,157,0,6,157,2,7,158,0,1,158,1,2,220,2,4,234,0,2,234,2,1,236,0,2,310,3,13,310,4,3,
/* out0389_em-eta9-phi19*/	10,91,2,4,157,0,10,220,0,2,220,1,9,220,2,8,233,2,1,234,2,5,236,0,3,236,1,11,310,3,3,
/* out0390_em-eta10-phi19*/	10,91,1,8,91,2,2,156,0,1,219,0,2,219,2,7,220,0,1,220,1,6,233,1,6,233,2,9,236,1,2,
/* out0391_em-eta11-phi19*/	11,35,2,13,35,3,10,35,4,1,35,5,1,91,1,4,156,0,1,219,0,11,219,1,1,219,2,1,232,2,4,233,1,9,
/* out0392_em-eta12-phi19*/	13,34,2,13,34,3,1,35,0,6,35,3,2,35,4,13,176,1,3,176,2,4,218,0,1,219,0,2,219,1,1,232,0,5,232,1,1,232,2,6,
/* out0393_em-eta13-phi19*/	9,34,1,12,34,2,3,35,0,3,35,1,9,176,1,6,218,0,3,227,2,1,232,0,6,232,1,2,
/* out0394_em-eta14-phi19*/	11,32,3,9,33,3,4,34,1,1,35,1,1,44,5,7,45,5,3,175,2,7,227,1,4,227,2,1,231,0,3,231,2,1,
/* out0395_em-eta15-phi19*/	10,32,0,10,32,3,4,44,4,4,44,5,1,175,0,2,175,1,2,175,2,2,226,2,1,227,1,3,231,0,3,
/* out0396_em-eta16-phi19*/	7,32,0,5,43,2,10,43,5,2,175,0,2,175,1,4,226,1,4,226,2,1,
/* out0397_em-eta17-phi19*/	6,43,0,1,43,4,6,43,5,6,175,1,1,226,0,2,226,1,3,
/* out0398_em-eta18-phi19*/	4,42,5,2,43,0,9,43,1,7,226,0,4,
/* out0399_em-eta19-phi19*/	3,42,4,3,43,0,1,43,1,6,
/* out0400_em-eta0-phi20*/	1,317,0,4,
/* out0401_em-eta1-phi20*/	2,317,0,12,317,1,6,
/* out0402_em-eta2-phi20*/	8,144,2,1,155,0,8,155,1,1,155,2,11,162,1,6,162,2,4,316,0,7,317,1,10,
/* out0403_em-eta3-phi20*/	9,154,0,6,154,2,2,155,0,8,155,1,5,161,1,11,161,2,11,162,1,1,316,0,9,316,1,9,
/* out0404_em-eta4-phi20*/	7,154,0,6,160,0,5,160,1,7,160,2,16,161,1,4,315,0,10,316,1,7,
/* out0405_em-eta5-phi20*/	8,94,1,2,94,2,1,159,0,6,159,2,10,160,0,4,160,1,8,315,0,6,315,1,11,
/* out0406_em-eta6-phi20*/	8,93,1,2,93,2,6,158,0,1,158,2,2,159,0,10,159,1,5,314,0,12,315,1,5,
/* out0407_em-eta7-phi20*/	5,92,2,4,93,1,8,158,0,9,314,0,4,314,1,13,
/* out0408_em-eta8-phi20*/	9,92,0,2,92,1,7,92,2,9,178,2,2,220,2,2,234,0,10,234,1,1,314,1,3,314,2,13,
/* out0409_em-eta9-phi20*/	10,91,0,1,91,2,7,92,1,7,178,1,5,220,0,10,220,2,2,234,0,3,234,1,7,234,2,10,314,2,3,
/* out0410_em-eta10-phi20*/	10,91,0,8,91,1,2,91,2,3,177,1,3,177,2,9,220,0,3,229,1,1,229,2,1,233,0,8,233,2,6,
/* out0411_em-eta11-phi20*/	12,34,3,2,35,3,4,46,5,4,47,5,7,91,0,3,91,1,2,176,2,2,177,1,10,219,0,1,228,2,4,233,0,8,233,1,1,
/* out0412_em-eta12-phi20*/	9,34,0,8,34,3,13,46,4,5,46,5,7,176,0,1,176,2,9,228,1,7,228,2,1,232,0,3,
/* out0413_em-eta13-phi20*/	10,34,0,8,34,1,3,45,2,10,45,5,6,46,4,1,176,0,4,176,1,5,227,2,6,228,1,2,232,0,2,
/* out0414_em-eta14-phi20*/	11,44,5,5,45,0,5,45,4,6,45,5,7,175,0,2,175,2,3,176,0,1,176,1,2,227,0,1,227,1,3,227,2,4,
/* out0415_em-eta15-phi20*/	6,44,4,9,44,5,3,45,0,4,45,1,4,175,0,6,227,1,6,
/* out0416_em-eta16-phi20*/	7,43,2,6,43,3,6,44,4,3,45,1,2,170,1,2,175,0,4,226,2,6,
/* out0417_em-eta17-phi20*/	6,42,2,2,43,3,3,43,4,9,170,1,3,226,0,3,226,2,3,
/* out0418_em-eta18-phi20*/	5,42,1,3,42,2,8,43,0,3,43,4,1,226,0,3,
/* out0419_em-eta19-phi20*/	4,42,1,4,42,2,2,43,0,2,43,1,3,
/* out0420_em-eta0-phi21*/	1,317,3,4,
/* out0421_em-eta1-phi21*/	2,317,2,6,317,3,12,
/* out0422_em-eta2-phi21*/	8,96,2,2,97,0,2,97,1,8,162,0,14,162,1,5,162,2,12,316,3,7,317,2,10,
/* out0423_em-eta3-phi21*/	9,95,2,3,96,1,12,96,2,8,161,0,13,161,2,5,162,0,2,162,1,4,316,2,9,316,3,9,
/* out0424_em-eta4-phi21*/	8,95,0,2,95,1,15,95,2,11,160,0,6,161,0,3,161,1,1,315,3,10,316,2,7,
/* out0425_em-eta5-phi21*/	7,94,0,7,94,1,7,94,2,15,95,1,1,160,0,1,315,2,11,315,3,6,
/* out0426_em-eta6-phi21*/	8,93,0,5,93,2,10,94,0,2,94,1,7,106,1,1,106,2,1,314,5,12,315,2,5,
/* out0427_em-eta7-phi21*/	6,92,2,1,93,0,10,93,1,6,105,2,3,314,4,13,314,5,4,
/* out0428_em-eta8-phi21*/	12,92,0,10,92,2,2,104,2,1,105,1,5,178,0,1,178,2,12,230,0,3,230,1,5,234,0,1,234,1,3,314,3,13,314,4,3,
/* out0429_em-eta9-phi21*/	11,91,0,1,92,0,4,104,1,3,104,2,7,178,0,7,178,1,10,178,2,2,229,2,8,230,1,7,234,1,5,314,3,3,
/* out0430_em-eta10-phi21*/	10,47,2,5,91,0,3,104,1,8,173,1,1,177,0,7,177,2,7,178,1,1,229,0,1,229,1,11,229,2,4,
/* out0431_em-eta11-phi21*/	12,46,5,1,47,0,1,47,2,11,47,3,5,47,4,14,47,5,9,172,2,2,177,0,8,177,1,3,228,0,1,228,2,9,229,1,3,
/* out0432_em-eta12-phi21*/	12,46,2,2,46,4,6,46,5,4,47,0,15,47,1,7,172,1,4,172,2,1,176,0,4,176,2,1,228,0,5,228,1,4,228,2,2,
/* out0433_em-eta13-phi21*/	12,45,2,6,45,3,13,45,4,1,46,4,4,47,1,5,171,2,3,172,1,1,176,0,6,227,0,1,227,2,3,228,0,1,228,1,3,
/* out0434_em-eta14-phi21*/	9,44,2,10,44,3,1,45,0,2,45,3,1,45,4,9,171,1,3,171,2,4,227,0,7,227,2,1,
/* out0435_em-eta15-phi21*/	7,44,1,6,44,2,5,45,0,5,45,1,4,171,1,6,222,2,1,227,0,5,
/* out0436_em-eta16-phi21*/	10,42,3,2,43,3,5,44,1,3,45,1,6,170,1,3,170,2,3,171,1,1,222,1,2,222,2,1,226,2,2,
/* out0437_em-eta17-phi21*/	7,42,2,1,42,3,11,43,3,2,170,1,5,222,1,2,226,0,1,226,2,3,
/* out0438_em-eta18-phi21*/	5,42,0,5,42,1,2,42,2,3,42,3,2,226,0,1,
/* out0439_em-eta19-phi21*/	2,42,0,2,42,1,7,
/* out0440_em-eta0-phi22*/	1,321,0,4,
/* out0441_em-eta1-phi22*/	2,321,0,12,321,1,6,
/* out0442_em-eta2-phi22*/	7,96,2,2,97,0,14,97,1,8,109,1,1,109,2,10,320,0,7,321,1,10,
/* out0443_em-eta3-phi22*/	9,95,2,1,96,0,16,96,1,4,96,2,4,108,1,1,108,2,12,109,1,10,320,0,9,320,1,9,
/* out0444_em-eta4-phi22*/	6,95,0,14,95,2,1,107,2,10,108,1,13,319,0,10,320,1,7,
/* out0445_em-eta5-phi22*/	7,94,0,6,106,2,4,107,0,2,107,1,15,107,2,4,319,0,6,319,1,11,
/* out0446_em-eta6-phi22*/	6,94,0,1,106,0,4,106,1,10,106,2,11,318,0,12,319,1,5,
/* out0447_em-eta7-phi22*/	7,93,0,1,105,0,3,105,2,12,106,0,1,106,1,5,318,0,4,318,1,13,
/* out0448_em-eta8-phi22*/	10,104,2,1,105,0,6,105,1,11,105,2,1,174,0,3,174,1,7,178,0,2,230,0,7,318,1,3,318,2,13,
/* out0449_em-eta9-phi22*/	12,104,0,7,104,2,7,173,2,9,174,1,6,178,0,6,225,1,3,225,2,4,229,0,2,229,2,3,230,0,6,230,1,4,318,2,3,
/* out0450_em-eta10-phi22*/	8,47,3,1,104,0,6,104,1,5,173,1,11,173,2,4,224,2,2,225,1,2,229,0,12,
/* out0451_em-eta11-phi22*/	13,46,0,3,46,2,5,46,3,15,47,3,10,47,4,2,172,2,9,173,1,2,177,0,1,224,1,5,224,2,4,228,0,2,229,0,1,229,1,1,
/* out0452_em-eta12-phi22*/	11,46,0,9,46,1,12,46,2,9,46,3,1,47,1,1,172,0,2,172,1,6,172,2,2,223,2,3,224,1,3,228,0,6,
/* out0453_em-eta13-phi22*/	9,44,3,5,45,3,2,46,1,4,47,1,3,171,2,5,172,1,4,223,1,3,223,2,6,228,0,1,
/* out0454_em-eta14-phi22*/	8,44,0,9,44,2,1,44,3,10,171,0,3,171,1,1,171,2,4,223,1,6,227,0,1,
/* out0455_em-eta15-phi22*/	6,44,0,7,44,1,6,171,0,2,171,1,4,222,2,6,227,0,1,
/* out0456_em-eta16-phi22*/	5,44,1,1,170,2,5,171,1,1,222,1,3,222,2,3,
/* out0457_em-eta17-phi22*/	5,42,0,1,42,3,1,170,1,2,170,2,4,222,1,5,
/* out0458_em-eta18-phi22*/	2,42,0,6,222,1,1,
/* out0459_em-eta19-phi22*/	1,42,0,2,
/* out0460_em-eta0-phi23*/	1,321,3,4,
/* out0461_em-eta1-phi23*/	2,321,2,6,321,3,12,
/* out0462_em-eta2-phi23*/	4,109,0,8,109,2,6,320,3,7,321,2,10,
/* out0463_em-eta3-phi23*/	6,108,0,7,108,2,4,109,0,8,109,1,5,320,2,9,320,3,9,
/* out0464_em-eta4-phi23*/	6,107,0,3,107,2,2,108,0,9,108,1,2,319,3,10,320,2,7,
/* out0465_em-eta5-phi23*/	4,107,0,11,107,1,1,319,2,11,319,3,6,
/* out0466_em-eta6-phi23*/	3,106,0,10,318,5,12,319,2,5,
/* out0467_em-eta7-phi23*/	4,105,0,3,106,0,1,318,4,13,318,5,4,
/* out0468_em-eta8-phi23*/	6,105,0,4,174,0,9,225,0,7,225,2,3,318,3,13,318,4,3,
/* out0469_em-eta9-phi23*/	9,104,0,2,173,0,3,173,2,3,174,0,4,174,1,3,225,0,7,225,1,4,225,2,9,318,3,3,
/* out0470_em-eta10-phi23*/	7,104,0,1,173,0,12,173,1,1,224,0,7,224,2,6,225,0,2,225,1,7,
/* out0471_em-eta11-phi23*/	8,46,0,1,172,0,4,172,2,2,173,0,1,173,1,1,224,0,7,224,1,3,224,2,4,
/* out0472_em-eta12-phi23*/	6,46,0,3,172,0,9,223,0,1,223,2,4,224,0,2,224,1,5,
/* out0473_em-eta13-phi23*/	6,171,0,1,172,0,1,172,1,1,223,0,6,223,1,1,223,2,3,
/* out0474_em-eta14-phi23*/	3,171,0,6,223,0,3,223,1,5,
/* out0475_em-eta15-phi23*/	5,171,0,4,222,0,2,222,2,4,223,0,6,223,1,1,
/* out0476_em-eta16-phi23*/	3,170,2,1,222,0,5,222,2,1,
/* out0477_em-eta17-phi23*/	3,170,2,3,222,0,3,222,1,2,
/* out0478_em-eta18-phi23*/	3,170,1,1,222,0,6,222,1,1,
/* out0479_em-eta19-phi23*/	0
};