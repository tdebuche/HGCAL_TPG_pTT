parameter integer matrixH [0:2382] = {
/* num inputs = 156(in0-in155) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 5 */
//* total number of input in adders 951 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	1, 133, 1, 
/* out0002_had-eta2-phi0*/	2, 132, 1, 133, 7, 
/* out0003_had-eta3-phi0*/	1, 132, 4, 
/* out0004_had-eta4-phi0*/	1, 132, 3, 
/* out0005_had-eta5-phi0*/	2, 93, 1, 94, 11, 
/* out0006_had-eta6-phi0*/	1, 93, 8, 
/* out0007_had-eta7-phi0*/	2, 92, 4, 93, 1, 
/* out0008_had-eta8-phi0*/	2, 91, 1, 92, 4, 
/* out0009_had-eta9-phi0*/	1, 91, 4, 
/* out0010_had-eta10-phi0*/	2, 90, 1, 91, 2, 
/* out0011_had-eta11-phi0*/	2, 90, 3, 127, 5, 
/* out0012_had-eta12-phi0*/	3, 90, 1, 126, 2, 127, 1, 
/* out0013_had-eta13-phi0*/	2, 89, 2, 126, 3, 
/* out0014_had-eta14-phi0*/	3, 89, 2, 125, 1, 126, 1, 
/* out0015_had-eta15-phi0*/	1, 125, 2, 
/* out0016_had-eta16-phi0*/	2, 88, 1, 125, 1, 
/* out0017_had-eta17-phi0*/	1, 88, 1, 
/* out0018_had-eta18-phi0*/	2, 88, 1, 124, 2, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	1, 133, 1, 
/* out0022_had-eta2-phi1*/	2, 132, 1, 133, 7, 
/* out0023_had-eta3-phi1*/	1, 132, 4, 
/* out0024_had-eta4-phi1*/	1, 132, 3, 
/* out0025_had-eta5-phi1*/	2, 87, 7, 94, 5, 
/* out0026_had-eta6-phi1*/	3, 86, 2, 87, 2, 93, 5, 
/* out0027_had-eta7-phi1*/	3, 86, 3, 92, 4, 93, 1, 
/* out0028_had-eta8-phi1*/	3, 85, 2, 91, 1, 92, 4, 
/* out0029_had-eta9-phi1*/	1, 91, 5, 
/* out0030_had-eta10-phi1*/	2, 90, 1, 91, 3, 
/* out0031_had-eta11-phi1*/	2, 90, 4, 127, 8, 
/* out0032_had-eta12-phi1*/	4, 89, 1, 90, 3, 126, 3, 127, 2, 
/* out0033_had-eta13-phi1*/	2, 89, 3, 126, 3, 
/* out0034_had-eta14-phi1*/	3, 89, 2, 125, 2, 126, 1, 
/* out0035_had-eta15-phi1*/	3, 88, 1, 89, 1, 125, 2, 
/* out0036_had-eta16-phi1*/	2, 88, 2, 125, 2, 
/* out0037_had-eta17-phi1*/	3, 88, 1, 124, 3, 125, 1, 
/* out0038_had-eta18-phi1*/	2, 88, 1, 124, 3, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	1, 135, 1, 
/* out0042_had-eta2-phi2*/	2, 134, 1, 135, 7, 
/* out0043_had-eta3-phi2*/	1, 134, 4, 
/* out0044_had-eta4-phi2*/	1, 134, 3, 
/* out0045_had-eta5-phi2*/	2, 81, 2, 87, 5, 
/* out0046_had-eta6-phi2*/	3, 81, 3, 86, 5, 87, 2, 
/* out0047_had-eta7-phi2*/	3, 80, 1, 85, 2, 86, 6, 
/* out0048_had-eta8-phi2*/	1, 85, 7, 
/* out0049_had-eta9-phi2*/	2, 84, 3, 85, 3, 
/* out0050_had-eta10-phi2*/	1, 84, 5, 
/* out0051_had-eta11-phi2*/	4, 83, 1, 84, 1, 90, 2, 122, 5, 
/* out0052_had-eta12-phi2*/	4, 83, 2, 90, 1, 122, 4, 126, 1, 
/* out0053_had-eta13-phi2*/	4, 83, 1, 89, 2, 121, 2, 126, 2, 
/* out0054_had-eta14-phi2*/	3, 89, 2, 121, 2, 125, 1, 
/* out0055_had-eta15-phi2*/	3, 88, 1, 89, 1, 125, 2, 
/* out0056_had-eta16-phi2*/	2, 88, 2, 125, 2, 
/* out0057_had-eta17-phi2*/	2, 88, 1, 124, 3, 
/* out0058_had-eta18-phi2*/	2, 88, 1, 124, 2, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 135, 1, 
/* out0062_had-eta2-phi3*/	2, 134, 1, 135, 7, 
/* out0063_had-eta3-phi3*/	1, 134, 4, 
/* out0064_had-eta4-phi3*/	1, 134, 3, 
/* out0065_had-eta5-phi3*/	2, 76, 8, 81, 4, 
/* out0066_had-eta6-phi3*/	3, 75, 1, 80, 2, 81, 7, 
/* out0067_had-eta7-phi3*/	1, 80, 8, 
/* out0068_had-eta8-phi3*/	3, 79, 3, 80, 2, 85, 2, 
/* out0069_had-eta9-phi3*/	2, 79, 3, 84, 2, 
/* out0070_had-eta10-phi3*/	1, 84, 4, 
/* out0071_had-eta11-phi3*/	3, 83, 3, 84, 1, 122, 4, 
/* out0072_had-eta12-phi3*/	3, 83, 3, 121, 1, 122, 3, 
/* out0073_had-eta13-phi3*/	3, 82, 1, 83, 2, 121, 3, 
/* out0074_had-eta14-phi3*/	2, 82, 2, 121, 3, 
/* out0075_had-eta15-phi3*/	3, 82, 2, 120, 2, 121, 1, 
/* out0076_had-eta16-phi3*/	2, 88, 1, 120, 2, 
/* out0077_had-eta17-phi3*/	3, 88, 1, 120, 1, 124, 1, 
/* out0078_had-eta18-phi3*/	2, 88, 1, 124, 2, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 137, 1, 
/* out0082_had-eta2-phi4*/	2, 136, 1, 137, 7, 
/* out0083_had-eta3-phi4*/	1, 136, 4, 
/* out0084_had-eta4-phi4*/	1, 136, 3, 
/* out0085_had-eta5-phi4*/	3, 75, 3, 76, 8, 77, 3, 
/* out0086_had-eta6-phi4*/	1, 75, 9, 
/* out0087_had-eta7-phi4*/	3, 74, 4, 75, 1, 80, 3, 
/* out0088_had-eta8-phi4*/	2, 74, 1, 79, 5, 
/* out0089_had-eta9-phi4*/	2, 78, 1, 79, 5, 
/* out0090_had-eta10-phi4*/	1, 78, 5, 
/* out0091_had-eta11-phi4*/	3, 78, 3, 83, 1, 123, 3, 
/* out0092_had-eta12-phi4*/	3, 63, 1, 83, 2, 123, 4, 
/* out0093_had-eta13-phi4*/	4, 82, 2, 83, 1, 121, 2, 123, 1, 
/* out0094_had-eta14-phi4*/	3, 82, 2, 116, 1, 121, 2, 
/* out0095_had-eta15-phi4*/	2, 82, 2, 120, 3, 
/* out0096_had-eta16-phi4*/	3, 49, 1, 82, 1, 120, 2, 
/* out0097_had-eta17-phi4*/	2, 49, 1, 120, 2, 
/* out0098_had-eta18-phi4*/	1, 49, 1, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 137, 1, 
/* out0102_had-eta2-phi5*/	2, 136, 1, 137, 7, 
/* out0103_had-eta3-phi5*/	1, 136, 4, 
/* out0104_had-eta4-phi5*/	1, 136, 3, 
/* out0105_had-eta5-phi5*/	2, 70, 1, 77, 13, 
/* out0106_had-eta6-phi5*/	3, 70, 6, 74, 1, 75, 2, 
/* out0107_had-eta7-phi5*/	1, 74, 7, 
/* out0108_had-eta8-phi5*/	2, 68, 3, 74, 3, 
/* out0109_had-eta9-phi5*/	2, 68, 4, 78, 1, 
/* out0110_had-eta10-phi5*/	1, 78, 4, 
/* out0111_had-eta11-phi5*/	3, 63, 2, 78, 2, 123, 3, 
/* out0112_had-eta12-phi5*/	2, 63, 3, 123, 4, 
/* out0113_had-eta13-phi5*/	3, 63, 2, 116, 3, 123, 1, 
/* out0114_had-eta14-phi5*/	2, 82, 2, 116, 3, 
/* out0115_had-eta15-phi5*/	3, 82, 2, 116, 1, 120, 1, 
/* out0116_had-eta16-phi5*/	2, 49, 2, 120, 2, 
/* out0117_had-eta17-phi5*/	2, 49, 2, 120, 1, 
/* out0118_had-eta18-phi5*/	1, 49, 1, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 139, 1, 
/* out0122_had-eta2-phi6*/	2, 138, 1, 139, 7, 
/* out0123_had-eta3-phi6*/	1, 138, 4, 
/* out0124_had-eta4-phi6*/	1, 138, 3, 
/* out0125_had-eta5-phi6*/	2, 70, 1, 72, 13, 
/* out0126_had-eta6-phi6*/	3, 69, 1, 70, 7, 71, 2, 
/* out0127_had-eta7-phi6*/	2, 69, 7, 70, 1, 
/* out0128_had-eta8-phi6*/	2, 68, 4, 69, 3, 
/* out0129_had-eta9-phi6*/	2, 64, 1, 68, 5, 
/* out0130_had-eta10-phi6*/	1, 64, 4, 
/* out0131_had-eta11-phi6*/	3, 63, 2, 64, 2, 118, 3, 
/* out0132_had-eta12-phi6*/	2, 63, 3, 118, 4, 
/* out0133_had-eta13-phi6*/	3, 63, 2, 116, 3, 118, 1, 
/* out0134_had-eta14-phi6*/	2, 50, 2, 116, 3, 
/* out0135_had-eta15-phi6*/	3, 50, 2, 115, 1, 116, 1, 
/* out0136_had-eta16-phi6*/	2, 49, 2, 115, 2, 
/* out0137_had-eta17-phi6*/	2, 49, 2, 115, 1, 
/* out0138_had-eta18-phi6*/	1, 49, 1, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 139, 1, 
/* out0142_had-eta2-phi7*/	2, 138, 1, 139, 7, 
/* out0143_had-eta3-phi7*/	1, 138, 4, 
/* out0144_had-eta4-phi7*/	1, 138, 3, 
/* out0145_had-eta5-phi7*/	3, 71, 3, 72, 3, 73, 8, 
/* out0146_had-eta6-phi7*/	1, 71, 9, 
/* out0147_had-eta7-phi7*/	3, 66, 3, 69, 4, 71, 1, 
/* out0148_had-eta8-phi7*/	2, 65, 5, 69, 1, 
/* out0149_had-eta9-phi7*/	2, 64, 1, 65, 5, 
/* out0150_had-eta10-phi7*/	1, 64, 5, 
/* out0151_had-eta11-phi7*/	3, 51, 1, 64, 3, 118, 3, 
/* out0152_had-eta12-phi7*/	3, 51, 2, 63, 1, 118, 4, 
/* out0153_had-eta13-phi7*/	4, 50, 2, 51, 1, 117, 2, 118, 1, 
/* out0154_had-eta14-phi7*/	3, 50, 2, 116, 1, 117, 2, 
/* out0155_had-eta15-phi7*/	2, 50, 2, 115, 3, 
/* out0156_had-eta16-phi7*/	3, 49, 1, 50, 1, 115, 2, 
/* out0157_had-eta17-phi7*/	2, 49, 1, 115, 2, 
/* out0158_had-eta18-phi7*/	1, 49, 1, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 141, 1, 
/* out0162_had-eta2-phi8*/	2, 140, 1, 141, 7, 
/* out0163_had-eta3-phi8*/	1, 140, 4, 
/* out0164_had-eta4-phi8*/	1, 140, 3, 
/* out0165_had-eta5-phi8*/	2, 67, 4, 73, 8, 
/* out0166_had-eta6-phi8*/	3, 66, 2, 67, 7, 71, 1, 
/* out0167_had-eta7-phi8*/	1, 66, 8, 
/* out0168_had-eta8-phi8*/	3, 53, 2, 65, 3, 66, 2, 
/* out0169_had-eta9-phi8*/	2, 52, 2, 65, 3, 
/* out0170_had-eta10-phi8*/	1, 52, 4, 
/* out0171_had-eta11-phi8*/	3, 51, 3, 52, 1, 119, 4, 
/* out0172_had-eta12-phi8*/	3, 51, 3, 117, 1, 119, 3, 
/* out0173_had-eta13-phi8*/	3, 50, 1, 51, 2, 117, 3, 
/* out0174_had-eta14-phi8*/	2, 50, 2, 117, 3, 
/* out0175_had-eta15-phi8*/	3, 50, 2, 115, 2, 117, 1, 
/* out0176_had-eta16-phi8*/	2, 56, 1, 115, 2, 
/* out0177_had-eta17-phi8*/	3, 56, 1, 111, 1, 115, 1, 
/* out0178_had-eta18-phi8*/	2, 56, 1, 111, 2, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 141, 1, 
/* out0182_had-eta2-phi9*/	2, 140, 1, 141, 7, 
/* out0183_had-eta3-phi9*/	1, 140, 4, 
/* out0184_had-eta4-phi9*/	1, 140, 3, 
/* out0185_had-eta5-phi9*/	2, 55, 5, 67, 2, 
/* out0186_had-eta6-phi9*/	3, 54, 5, 55, 2, 67, 3, 
/* out0187_had-eta7-phi9*/	3, 53, 2, 54, 6, 66, 1, 
/* out0188_had-eta8-phi9*/	1, 53, 7, 
/* out0189_had-eta9-phi9*/	2, 52, 3, 53, 3, 
/* out0190_had-eta10-phi9*/	1, 52, 5, 
/* out0191_had-eta11-phi9*/	4, 51, 1, 52, 1, 58, 2, 119, 5, 
/* out0192_had-eta12-phi9*/	4, 51, 2, 58, 1, 113, 1, 119, 4, 
/* out0193_had-eta13-phi9*/	4, 51, 1, 57, 2, 113, 2, 117, 2, 
/* out0194_had-eta14-phi9*/	3, 57, 2, 112, 1, 117, 2, 
/* out0195_had-eta15-phi9*/	3, 56, 1, 57, 1, 112, 2, 
/* out0196_had-eta16-phi9*/	2, 56, 2, 112, 2, 
/* out0197_had-eta17-phi9*/	2, 56, 1, 111, 3, 
/* out0198_had-eta18-phi9*/	2, 56, 1, 111, 2, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 143, 1, 
/* out0202_had-eta2-phi10*/	2, 142, 1, 143, 7, 
/* out0203_had-eta3-phi10*/	1, 142, 4, 
/* out0204_had-eta4-phi10*/	1, 142, 3, 
/* out0205_had-eta5-phi10*/	2, 55, 7, 62, 5, 
/* out0206_had-eta6-phi10*/	3, 54, 2, 55, 2, 61, 5, 
/* out0207_had-eta7-phi10*/	3, 54, 3, 60, 4, 61, 1, 
/* out0208_had-eta8-phi10*/	3, 53, 2, 59, 1, 60, 4, 
/* out0209_had-eta9-phi10*/	1, 59, 5, 
/* out0210_had-eta10-phi10*/	2, 58, 1, 59, 3, 
/* out0211_had-eta11-phi10*/	2, 58, 4, 114, 8, 
/* out0212_had-eta12-phi10*/	4, 57, 1, 58, 3, 113, 3, 114, 2, 
/* out0213_had-eta13-phi10*/	2, 57, 3, 113, 3, 
/* out0214_had-eta14-phi10*/	3, 57, 2, 112, 2, 113, 1, 
/* out0215_had-eta15-phi10*/	3, 56, 1, 57, 1, 112, 2, 
/* out0216_had-eta16-phi10*/	2, 56, 2, 112, 2, 
/* out0217_had-eta17-phi10*/	3, 56, 1, 111, 3, 112, 1, 
/* out0218_had-eta18-phi10*/	2, 56, 1, 111, 3, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 143, 1, 
/* out0222_had-eta2-phi11*/	2, 142, 1, 143, 7, 
/* out0223_had-eta3-phi11*/	1, 142, 4, 
/* out0224_had-eta4-phi11*/	1, 142, 3, 
/* out0225_had-eta5-phi11*/	3, 48, 2, 61, 1, 62, 11, 
/* out0226_had-eta6-phi11*/	3, 47, 1, 48, 1, 61, 8, 
/* out0227_had-eta7-phi11*/	3, 47, 2, 60, 4, 61, 1, 
/* out0228_had-eta8-phi11*/	3, 46, 2, 59, 1, 60, 4, 
/* out0229_had-eta9-phi11*/	2, 46, 1, 59, 4, 
/* out0230_had-eta10-phi11*/	3, 45, 2, 58, 1, 59, 2, 
/* out0231_had-eta11-phi11*/	4, 45, 1, 58, 3, 110, 1, 114, 5, 
/* out0232_had-eta12-phi11*/	5, 44, 1, 58, 1, 110, 2, 113, 2, 114, 1, 
/* out0233_had-eta13-phi11*/	3, 44, 1, 57, 2, 113, 3, 
/* out0234_had-eta14-phi11*/	4, 57, 2, 109, 2, 112, 1, 113, 1, 
/* out0235_had-eta15-phi11*/	3, 43, 1, 109, 1, 112, 2, 
/* out0236_had-eta16-phi11*/	4, 43, 1, 56, 1, 108, 1, 112, 1, 
/* out0237_had-eta17-phi11*/	2, 56, 1, 108, 1, 
/* out0238_had-eta18-phi11*/	4, 42, 1, 56, 1, 108, 1, 111, 2, 
/* out0239_had-eta19-phi11*/	1, 42, 1, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 145, 1, 
/* out0242_had-eta2-phi12*/	2, 144, 1, 145, 7, 
/* out0243_had-eta3-phi12*/	1, 144, 4, 
/* out0244_had-eta4-phi12*/	1, 144, 3, 
/* out0245_had-eta5-phi12*/	2, 41, 1, 48, 8, 
/* out0246_had-eta6-phi12*/	3, 40, 1, 47, 4, 48, 5, 
/* out0247_had-eta7-phi12*/	1, 47, 8, 
/* out0248_had-eta8-phi12*/	1, 46, 6, 
/* out0249_had-eta9-phi12*/	2, 45, 1, 46, 4, 
/* out0250_had-eta10-phi12*/	1, 45, 5, 
/* out0251_had-eta11-phi12*/	3, 44, 1, 45, 3, 110, 4, 
/* out0252_had-eta12-phi12*/	2, 44, 3, 110, 4, 
/* out0253_had-eta13-phi12*/	3, 44, 3, 109, 2, 110, 1, 
/* out0254_had-eta14-phi12*/	3, 43, 2, 44, 1, 109, 3, 
/* out0255_had-eta15-phi12*/	2, 43, 2, 109, 2, 
/* out0256_had-eta16-phi12*/	2, 43, 2, 108, 2, 
/* out0257_had-eta17-phi12*/	3, 42, 1, 43, 1, 108, 2, 
/* out0258_had-eta18-phi12*/	2, 42, 2, 108, 2, 
/* out0259_had-eta19-phi12*/	1, 42, 1, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 145, 1, 
/* out0262_had-eta2-phi13*/	2, 144, 1, 145, 7, 
/* out0263_had-eta3-phi13*/	1, 144, 4, 
/* out0264_had-eta4-phi13*/	1, 144, 3, 
/* out0265_had-eta5-phi13*/	2, 40, 2, 41, 14, 
/* out0266_had-eta6-phi13*/	1, 40, 9, 
/* out0267_had-eta7-phi13*/	3, 39, 6, 40, 1, 47, 1, 
/* out0268_had-eta8-phi13*/	3, 38, 1, 39, 4, 46, 2, 
/* out0269_had-eta9-phi13*/	2, 38, 4, 46, 1, 
/* out0270_had-eta10-phi13*/	3, 37, 1, 38, 1, 45, 3, 
/* out0271_had-eta11-phi13*/	5, 37, 2, 44, 1, 45, 1, 107, 5, 110, 1, 
/* out0272_had-eta12-phi13*/	4, 44, 3, 105, 1, 107, 1, 110, 3, 
/* out0273_had-eta13-phi13*/	3, 44, 2, 105, 2, 109, 1, 
/* out0274_had-eta14-phi13*/	2, 43, 2, 109, 3, 
/* out0275_had-eta15-phi13*/	3, 43, 2, 103, 1, 109, 2, 
/* out0276_had-eta16-phi13*/	2, 43, 1, 108, 2, 
/* out0277_had-eta17-phi13*/	2, 42, 2, 108, 2, 
/* out0278_had-eta18-phi13*/	2, 42, 2, 108, 1, 
/* out0279_had-eta19-phi13*/	1, 42, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 147, 1, 
/* out0282_had-eta2-phi14*/	2, 146, 1, 147, 7, 
/* out0283_had-eta3-phi14*/	1, 146, 4, 
/* out0284_had-eta4-phi14*/	1, 146, 3, 
/* out0285_had-eta5-phi14*/	2, 24, 10, 41, 1, 
/* out0286_had-eta6-phi14*/	3, 23, 5, 24, 2, 40, 3, 
/* out0287_had-eta7-phi14*/	3, 22, 1, 23, 3, 39, 4, 
/* out0288_had-eta8-phi14*/	3, 22, 2, 38, 2, 39, 2, 
/* out0289_had-eta9-phi14*/	1, 38, 5, 
/* out0290_had-eta10-phi14*/	2, 37, 2, 38, 2, 
/* out0291_had-eta11-phi14*/	2, 37, 4, 107, 9, 
/* out0292_had-eta12-phi14*/	3, 36, 1, 37, 2, 105, 4, 
/* out0293_had-eta13-phi14*/	2, 36, 3, 105, 4, 
/* out0294_had-eta14-phi14*/	3, 36, 2, 103, 2, 105, 1, 
/* out0295_had-eta15-phi14*/	2, 43, 1, 103, 2, 
/* out0296_had-eta16-phi14*/	4, 35, 1, 43, 1, 103, 1, 108, 1, 
/* out0297_had-eta17-phi14*/	4, 35, 1, 42, 1, 102, 1, 108, 1, 
/* out0298_had-eta18-phi14*/	2, 42, 2, 102, 1, 
/* out0299_had-eta19-phi14*/	1, 42, 1, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 147, 1, 
/* out0302_had-eta2-phi15*/	2, 146, 1, 147, 7, 
/* out0303_had-eta3-phi15*/	1, 146, 4, 
/* out0304_had-eta4-phi15*/	1, 146, 3, 
/* out0305_had-eta5-phi15*/	2, 24, 3, 28, 5, 
/* out0306_had-eta6-phi15*/	4, 23, 5, 24, 1, 26, 1, 28, 4, 
/* out0307_had-eta7-phi15*/	3, 22, 3, 23, 3, 26, 2, 
/* out0308_had-eta8-phi15*/	1, 22, 7, 
/* out0309_had-eta9-phi15*/	3, 21, 4, 22, 1, 38, 1, 
/* out0310_had-eta10-phi15*/	2, 21, 4, 37, 1, 
/* out0311_had-eta11-phi15*/	4, 20, 1, 37, 3, 106, 6, 107, 1, 
/* out0312_had-eta12-phi15*/	5, 20, 1, 36, 2, 37, 1, 105, 2, 106, 2, 
/* out0313_had-eta13-phi15*/	3, 36, 3, 104, 1, 105, 2, 
/* out0314_had-eta14-phi15*/	2, 36, 2, 103, 3, 
/* out0315_had-eta15-phi15*/	2, 35, 1, 103, 2, 
/* out0316_had-eta16-phi15*/	2, 35, 2, 103, 2, 
/* out0317_had-eta17-phi15*/	2, 35, 1, 102, 2, 
/* out0318_had-eta18-phi15*/	3, 35, 1, 42, 1, 102, 2, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 149, 1, 
/* out0322_had-eta2-phi16*/	2, 148, 1, 149, 7, 
/* out0323_had-eta3-phi16*/	1, 148, 4, 
/* out0324_had-eta4-phi16*/	1, 148, 3, 
/* out0325_had-eta5-phi16*/	2, 27, 2, 28, 4, 
/* out0326_had-eta6-phi16*/	3, 26, 5, 27, 2, 28, 3, 
/* out0327_had-eta7-phi16*/	2, 25, 1, 26, 7, 
/* out0328_had-eta8-phi16*/	2, 22, 2, 25, 5, 
/* out0329_had-eta9-phi16*/	2, 21, 4, 25, 1, 
/* out0330_had-eta10-phi16*/	2, 20, 1, 21, 4, 
/* out0331_had-eta11-phi16*/	2, 20, 4, 106, 5, 
/* out0332_had-eta12-phi16*/	3, 20, 3, 104, 2, 106, 3, 
/* out0333_had-eta13-phi16*/	3, 14, 1, 36, 2, 104, 4, 
/* out0334_had-eta14-phi16*/	4, 14, 1, 36, 1, 103, 1, 104, 2, 
/* out0335_had-eta15-phi16*/	3, 35, 2, 98, 1, 103, 1, 
/* out0336_had-eta16-phi16*/	4, 35, 2, 98, 1, 102, 1, 103, 1, 
/* out0337_had-eta17-phi16*/	2, 35, 1, 102, 2, 
/* out0338_had-eta18-phi16*/	2, 35, 1, 102, 2, 
/* out0339_had-eta19-phi16*/	1, 102, 1, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 149, 1, 
/* out0342_had-eta2-phi17*/	2, 148, 1, 149, 7, 
/* out0343_had-eta3-phi17*/	1, 148, 4, 
/* out0344_had-eta4-phi17*/	1, 148, 3, 
/* out0345_had-eta5-phi17*/	1, 27, 6, 
/* out0346_had-eta6-phi17*/	2, 27, 6, 33, 2, 
/* out0347_had-eta7-phi17*/	3, 25, 1, 26, 1, 33, 5, 
/* out0348_had-eta8-phi17*/	1, 25, 6, 
/* out0349_had-eta9-phi17*/	2, 25, 2, 29, 3, 
/* out0350_had-eta10-phi17*/	1, 29, 4, 
/* out0351_had-eta11-phi17*/	2, 20, 3, 101, 5, 
/* out0352_had-eta12-phi17*/	3, 20, 3, 101, 3, 104, 2, 
/* out0353_had-eta13-phi17*/	2, 14, 3, 104, 3, 
/* out0354_had-eta14-phi17*/	3, 14, 2, 98, 1, 104, 2, 
/* out0355_had-eta15-phi17*/	3, 14, 1, 35, 1, 98, 3, 
/* out0356_had-eta16-phi17*/	2, 35, 1, 98, 2, 
/* out0357_had-eta17-phi17*/	2, 35, 1, 102, 1, 
/* out0358_had-eta18-phi17*/	1, 102, 2, 
/* out0359_had-eta19-phi17*/	1, 102, 1, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 151, 1, 
/* out0362_had-eta2-phi18*/	2, 150, 1, 151, 7, 
/* out0363_had-eta3-phi18*/	1, 150, 4, 
/* out0364_had-eta4-phi18*/	1, 150, 3, 
/* out0365_had-eta5-phi18*/	1, 34, 6, 
/* out0366_had-eta6-phi18*/	2, 33, 3, 34, 6, 
/* out0367_had-eta7-phi18*/	3, 30, 1, 31, 1, 33, 6, 
/* out0368_had-eta8-phi18*/	1, 30, 6, 
/* out0369_had-eta9-phi18*/	2, 29, 4, 30, 2, 
/* out0370_had-eta10-phi18*/	1, 29, 4, 
/* out0371_had-eta11-phi18*/	3, 15, 3, 29, 1, 101, 5, 
/* out0372_had-eta12-phi18*/	3, 15, 3, 99, 2, 101, 3, 
/* out0373_had-eta13-phi18*/	2, 14, 3, 99, 3, 
/* out0374_had-eta14-phi18*/	3, 14, 2, 98, 1, 99, 2, 
/* out0375_had-eta15-phi18*/	3, 7, 1, 14, 1, 98, 3, 
/* out0376_had-eta16-phi18*/	2, 7, 1, 98, 2, 
/* out0377_had-eta17-phi18*/	2, 7, 1, 128, 1, 
/* out0378_had-eta18-phi18*/	1, 128, 2, 
/* out0379_had-eta19-phi18*/	1, 128, 1, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 151, 1, 
/* out0382_had-eta2-phi19*/	2, 150, 1, 151, 7, 
/* out0383_had-eta3-phi19*/	1, 150, 4, 
/* out0384_had-eta4-phi19*/	1, 150, 3, 
/* out0385_had-eta5-phi19*/	2, 32, 4, 34, 2, 
/* out0386_had-eta6-phi19*/	3, 31, 5, 32, 3, 34, 2, 
/* out0387_had-eta7-phi19*/	2, 30, 1, 31, 7, 
/* out0388_had-eta8-phi19*/	2, 17, 2, 30, 5, 
/* out0389_had-eta9-phi19*/	2, 16, 4, 30, 1, 
/* out0390_had-eta10-phi19*/	2, 15, 1, 16, 4, 
/* out0391_had-eta11-phi19*/	2, 15, 4, 100, 5, 
/* out0392_had-eta12-phi19*/	3, 15, 3, 99, 2, 100, 3, 
/* out0393_had-eta13-phi19*/	3, 8, 2, 14, 1, 99, 4, 
/* out0394_had-eta14-phi19*/	4, 8, 1, 14, 1, 99, 2, 129, 1, 
/* out0395_had-eta15-phi19*/	3, 7, 2, 98, 1, 129, 1, 
/* out0396_had-eta16-phi19*/	4, 7, 2, 98, 1, 128, 1, 129, 1, 
/* out0397_had-eta17-phi19*/	2, 7, 1, 128, 2, 
/* out0398_had-eta18-phi19*/	2, 7, 1, 128, 2, 
/* out0399_had-eta19-phi19*/	1, 128, 1, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 153, 1, 
/* out0402_had-eta2-phi20*/	2, 152, 1, 153, 7, 
/* out0403_had-eta3-phi20*/	1, 152, 4, 
/* out0404_had-eta4-phi20*/	1, 152, 3, 
/* out0405_had-eta5-phi20*/	2, 19, 3, 32, 5, 
/* out0406_had-eta6-phi20*/	4, 18, 5, 19, 1, 31, 1, 32, 4, 
/* out0407_had-eta7-phi20*/	3, 17, 3, 18, 3, 31, 2, 
/* out0408_had-eta8-phi20*/	1, 17, 7, 
/* out0409_had-eta9-phi20*/	3, 10, 1, 16, 4, 17, 1, 
/* out0410_had-eta10-phi20*/	2, 9, 1, 16, 4, 
/* out0411_had-eta11-phi20*/	4, 9, 3, 15, 1, 100, 6, 131, 1, 
/* out0412_had-eta12-phi20*/	5, 8, 2, 9, 1, 15, 1, 100, 2, 130, 2, 
/* out0413_had-eta13-phi20*/	3, 8, 3, 99, 1, 130, 2, 
/* out0414_had-eta14-phi20*/	2, 8, 2, 129, 3, 
/* out0415_had-eta15-phi20*/	2, 7, 1, 129, 2, 
/* out0416_had-eta16-phi20*/	2, 7, 2, 129, 2, 
/* out0417_had-eta17-phi20*/	2, 7, 1, 128, 2, 
/* out0418_had-eta18-phi20*/	3, 0, 1, 7, 1, 128, 2, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 153, 1, 
/* out0422_had-eta2-phi21*/	2, 152, 1, 153, 7, 
/* out0423_had-eta3-phi21*/	1, 152, 4, 
/* out0424_had-eta4-phi21*/	1, 152, 3, 
/* out0425_had-eta5-phi21*/	2, 13, 1, 19, 10, 
/* out0426_had-eta6-phi21*/	3, 12, 3, 18, 5, 19, 2, 
/* out0427_had-eta7-phi21*/	3, 11, 4, 17, 1, 18, 3, 
/* out0428_had-eta8-phi21*/	3, 10, 2, 11, 2, 17, 2, 
/* out0429_had-eta9-phi21*/	1, 10, 5, 
/* out0430_had-eta10-phi21*/	2, 9, 2, 10, 2, 
/* out0431_had-eta11-phi21*/	2, 9, 4, 131, 9, 
/* out0432_had-eta12-phi21*/	3, 8, 1, 9, 2, 130, 4, 
/* out0433_had-eta13-phi21*/	2, 8, 3, 130, 4, 
/* out0434_had-eta14-phi21*/	3, 8, 2, 129, 2, 130, 1, 
/* out0435_had-eta15-phi21*/	2, 1, 1, 129, 2, 
/* out0436_had-eta16-phi21*/	4, 1, 1, 7, 1, 95, 1, 129, 1, 
/* out0437_had-eta17-phi21*/	4, 0, 1, 7, 1, 95, 1, 128, 1, 
/* out0438_had-eta18-phi21*/	3, 0, 2, 95, 1, 128, 1, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 155, 1, 
/* out0442_had-eta2-phi22*/	2, 154, 1, 155, 7, 
/* out0443_had-eta3-phi22*/	1, 154, 4, 
/* out0444_had-eta4-phi22*/	1, 154, 3, 
/* out0445_had-eta5-phi22*/	3, 6, 1, 12, 2, 13, 14, 
/* out0446_had-eta6-phi22*/	1, 12, 9, 
/* out0447_had-eta7-phi22*/	3, 5, 2, 11, 6, 12, 1, 
/* out0448_had-eta8-phi22*/	3, 4, 2, 10, 1, 11, 4, 
/* out0449_had-eta9-phi22*/	3, 3, 1, 4, 1, 10, 4, 
/* out0450_had-eta10-phi22*/	3, 3, 3, 9, 1, 10, 1, 
/* out0451_had-eta11-phi22*/	5, 2, 1, 3, 2, 9, 2, 97, 2, 131, 5, 
/* out0452_had-eta12-phi22*/	4, 2, 3, 97, 3, 130, 1, 131, 1, 
/* out0453_had-eta13-phi22*/	3, 2, 3, 96, 2, 130, 2, 
/* out0454_had-eta14-phi22*/	2, 1, 2, 96, 3, 
/* out0455_had-eta15-phi22*/	4, 1, 2, 95, 1, 96, 2, 129, 1, 
/* out0456_had-eta16-phi22*/	2, 1, 2, 95, 2, 
/* out0457_had-eta17-phi22*/	3, 0, 2, 1, 1, 95, 2, 
/* out0458_had-eta18-phi22*/	2, 0, 3, 95, 2, 
/* out0459_had-eta19-phi22*/	1, 0, 1, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 155, 1, 
/* out0462_had-eta2-phi23*/	2, 154, 1, 155, 7, 
/* out0463_had-eta3-phi23*/	1, 154, 4, 
/* out0464_had-eta4-phi23*/	1, 154, 3, 
/* out0465_had-eta5-phi23*/	2, 6, 9, 13, 1, 
/* out0466_had-eta6-phi23*/	3, 5, 5, 6, 6, 12, 1, 
/* out0467_had-eta7-phi23*/	1, 5, 9, 
/* out0468_had-eta8-phi23*/	1, 4, 8, 
/* out0469_had-eta9-phi23*/	2, 3, 2, 4, 5, 
/* out0470_had-eta10-phi23*/	1, 3, 5, 
/* out0471_had-eta11-phi23*/	3, 2, 1, 3, 3, 97, 4, 
/* out0472_had-eta12-phi23*/	2, 2, 4, 97, 5, 
/* out0473_had-eta13-phi23*/	3, 2, 3, 96, 3, 97, 2, 
/* out0474_had-eta14-phi23*/	3, 1, 2, 2, 1, 96, 3, 
/* out0475_had-eta15-phi23*/	2, 1, 2, 96, 3, 
/* out0476_had-eta16-phi23*/	2, 1, 2, 95, 2, 
/* out0477_had-eta17-phi23*/	3, 0, 2, 1, 1, 95, 2, 
/* out0478_had-eta18-phi23*/	2, 0, 3, 95, 2, 
/* out0479_had-eta19-phi23*/	1, 0, 1, 
};