parameter integer matrixH [0:8939] = {
/* num inputs = 163(in0-in162) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 15 */
//* total number of input in adders 2819 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	2,82,1,4,82,2,7,
/* out0003_em-eta3-phi0*/	4,81,0,6,81,1,15,81,2,4,82,1,10,
/* out0004_em-eta4-phi0*/	4,63,0,4,63,1,3,81,0,10,81,2,7,
/* out0005_em-eta5-phi0*/	7,62,0,3,62,1,13,63,0,4,79,0,16,79,1,11,79,2,3,89,2,3,
/* out0006_em-eta6-phi0*/	9,42,0,1,62,0,13,62,2,5,68,0,10,68,1,4,79,1,4,79,2,13,80,0,1,80,2,1,
/* out0007_em-eta7-phi0*/	6,41,1,1,42,0,3,57,0,5,68,0,6,68,1,8,68,2,16,
/* out0008_em-eta8-phi0*/	5,41,0,6,41,1,9,57,0,11,57,1,6,57,2,3,
/* out0009_em-eta9-phi0*/	4,41,0,10,46,0,6,57,1,2,57,2,10,
/* out0010_em-eta10-phi0*/	3,46,0,7,46,1,3,46,2,7,
/* out0011_em-eta11-phi0*/	4,20,0,7,20,1,9,35,0,4,46,2,8,
/* out0012_em-eta12-phi0*/	8,20,0,9,20,1,1,20,2,9,20,3,12,21,4,1,35,0,8,35,1,1,35,2,1,
/* out0013_em-eta13-phi0*/	4,20,3,4,21,2,1,21,3,13,35,2,8,
/* out0014_em-eta14-phi0*/	2,24,0,8,35,2,4,
/* out0015_em-eta15-phi0*/	2,24,0,4,24,2,2,
/* out0016_em-eta16-phi0*/	2,1,1,2,24,2,5,
/* out0017_em-eta17-phi0*/	4,0,1,7,1,1,6,14,2,3,24,2,2,
/* out0018_em-eta18-phi0*/	3,0,0,4,0,1,8,14,2,5,
/* out0019_em-eta19-phi0*/	3,0,0,9,14,0,2,14,2,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	4,65,1,6,65,2,5,82,0,6,82,2,9,
/* out0023_em-eta3-phi1*/	8,64,0,15,64,1,7,64,2,3,65,1,5,81,1,1,81,2,3,82,0,10,82,1,2,
/* out0024_em-eta4-phi1*/	7,44,0,1,63,0,2,63,1,13,63,2,8,64,0,1,64,2,9,81,2,2,
/* out0025_em-eta5-phi1*/	11,43,0,10,62,1,3,62,2,3,63,0,6,63,2,8,79,1,1,80,0,7,80,1,1,89,1,14,89,2,13,90,0,1,
/* out0026_em-eta6-phi1*/	9,42,0,5,42,1,5,43,0,3,43,2,3,62,2,8,68,1,1,80,0,8,80,1,5,80,2,14,
/* out0027_em-eta7-phi1*/	8,42,0,7,42,1,3,42,2,11,68,1,3,69,0,15,69,1,1,69,2,3,80,2,1,
/* out0028_em-eta8-phi1*/	7,23,0,2,41,1,6,41,2,8,42,2,1,57,1,6,58,0,4,69,2,10,
/* out0029_em-eta9-phi1*/	8,22,1,5,41,2,8,46,0,3,46,1,1,57,1,2,57,2,3,58,0,7,58,2,5,
/* out0030_em-eta10-phi1*/	5,22,0,9,22,1,2,46,1,9,47,0,2,58,2,3,
/* out0031_em-eta11-phi1*/	12,20,1,6,20,2,1,20,4,3,21,0,1,21,1,16,22,0,3,35,0,1,35,1,1,46,1,3,46,2,1,47,0,4,47,2,2,
/* out0032_em-eta12-phi1*/	7,20,2,6,20,5,1,21,0,15,21,4,10,35,0,3,35,1,8,47,2,1,
/* out0033_em-eta13-phi1*/	8,2,0,1,21,2,14,21,3,3,21,4,5,21,5,5,35,1,5,35,2,2,36,0,1,
/* out0034_em-eta14-phi1*/	7,2,0,9,2,3,1,21,2,1,24,0,3,24,1,3,35,2,1,36,2,1,
/* out0035_em-eta15-phi1*/	4,2,3,5,24,0,1,24,1,5,24,2,1,
/* out0036_em-eta16-phi1*/	4,0,4,10,1,1,2,24,1,2,24,2,3,
/* out0037_em-eta17-phi1*/	5,0,2,1,1,0,7,1,1,6,14,2,3,24,2,2,
/* out0038_em-eta18-phi1*/	5,0,0,1,0,1,1,0,2,10,14,0,3,14,2,2,
/* out0039_em-eta19-phi1*/	4,0,0,2,0,2,1,0,3,6,14,0,2,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	5,46,0,1,46,1,9,65,0,11,65,1,1,65,2,11,
/* out0043_em-eta3-phi2*/	6,45,0,13,45,1,12,64,1,9,64,2,1,65,0,5,65,1,4,
/* out0044_em-eta4-phi2*/	5,44,0,14,44,1,11,44,2,6,45,0,2,64,2,3,
/* out0045_em-eta5-phi2*/	12,25,0,2,25,1,1,43,0,3,43,1,15,43,2,1,44,0,1,44,2,8,80,1,1,89,1,2,90,0,15,90,1,10,90,2,11,
/* out0046_em-eta6-phi2*/	9,24,0,3,24,1,6,42,1,3,43,1,1,43,2,12,80,1,9,81,0,14,81,2,2,90,2,4,
/* out0047_em-eta7-phi2*/	9,23,0,3,23,1,3,24,0,7,42,1,5,42,2,4,69,0,1,69,1,12,70,0,2,81,2,8,
/* out0048_em-eta8-phi2*/	9,23,0,11,23,1,3,23,2,3,58,0,3,58,1,3,69,1,3,69,2,3,70,0,4,70,2,3,
/* out0049_em-eta9-phi2*/	6,22,1,7,22,2,1,23,2,6,58,0,2,58,1,10,58,2,4,
/* out0050_em-eta10-phi2*/	7,22,0,2,22,1,2,22,2,8,47,0,7,47,1,2,58,1,1,58,2,4,
/* out0051_em-eta11-phi2*/	8,4,1,5,5,1,7,20,4,8,22,0,2,22,2,3,47,0,3,47,1,2,47,2,5,
/* out0052_em-eta12-phi2*/	8,4,0,6,4,1,6,20,4,5,20,5,15,21,5,2,35,1,1,36,0,3,47,2,6,
/* out0053_em-eta13-phi2*/	6,2,0,2,2,1,13,3,1,2,4,0,1,21,5,9,36,0,7,
/* out0054_em-eta14-phi2*/	6,2,0,4,2,1,3,2,2,12,2,3,4,24,1,1,36,2,6,
/* out0055_em-eta15-phi2*/	7,2,2,2,2,3,6,3,3,9,3,4,2,24,1,3,25,0,1,36,2,1,
/* out0056_em-eta16-phi2*/	5,0,4,6,0,5,6,3,3,4,24,1,2,25,0,3,
/* out0057_em-eta17-phi2*/	8,0,5,3,1,0,8,1,4,2,14,0,2,14,2,2,24,2,1,25,0,1,25,2,2,
/* out0058_em-eta18-phi2*/	5,0,2,2,1,0,1,1,3,3,1,4,8,14,0,4,
/* out0059_em-eta19-phi2*/	5,0,2,2,0,3,10,1,3,4,1,4,2,14,0,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	3,27,1,5,46,0,12,46,1,7,
/* out0063_em-eta3-phi3*/	6,26,1,6,27,0,12,27,1,5,45,1,4,45,2,15,46,0,3,
/* out0064_em-eta4-phi3*/	8,25,1,2,26,0,16,26,1,8,26,2,2,44,1,5,44,2,2,45,0,1,45,2,1,
/* out0065_em-eta5-phi3*/	6,25,0,9,25,1,13,25,2,8,90,1,6,91,0,15,91,2,2,
/* out0066_em-eta6-phi3*/	11,8,0,1,24,1,10,24,2,7,25,0,5,25,2,2,81,0,2,81,1,14,81,2,1,82,0,3,90,2,1,91,2,8,
/* out0067_em-eta7-phi3*/	11,7,0,1,7,1,3,23,1,2,24,0,6,24,2,8,70,0,7,70,1,5,81,1,2,81,2,5,82,0,2,82,2,2,
/* out0068_em-eta8-phi3*/	8,6,0,1,6,1,1,7,0,4,23,1,8,23,2,4,70,0,3,70,1,5,70,2,11,
/* out0069_em-eta9-phi3*/	6,6,0,10,22,2,1,23,2,3,58,1,2,59,0,13,70,2,2,
/* out0070_em-eta10-phi3*/	7,4,4,8,6,0,4,6,2,3,22,2,3,47,1,3,59,0,1,59,2,9,
/* out0071_em-eta11-phi3*/	9,4,1,1,4,2,2,4,4,8,4,5,4,5,0,14,5,1,9,5,4,1,47,1,8,48,0,3,
/* out0072_em-eta12-phi3*/	11,4,0,6,4,1,4,4,2,14,4,3,8,5,4,1,36,0,3,36,1,2,47,1,1,47,2,2,48,0,1,48,2,1,
/* out0073_em-eta13-phi3*/	7,2,4,6,3,0,1,3,1,14,4,0,3,4,3,4,36,0,2,36,1,5,
/* out0074_em-eta14-phi3*/	6,2,2,2,2,5,1,3,0,15,3,4,5,36,1,1,36,2,6,
/* out0075_em-eta15-phi3*/	6,3,2,5,3,3,3,3,4,9,3,5,3,25,0,4,36,2,1,
/* out0076_em-eta16-phi3*/	6,0,5,5,1,5,2,3,2,8,28,1,1,29,1,1,25,0,4,
/* out0077_em-eta17-phi3*/	4,0,5,2,1,4,1,1,5,11,25,2,4,
/* out0078_em-eta18-phi3*/	6,1,2,5,1,3,2,1,4,3,1,5,2,14,0,2,25,2,2,
/* out0079_em-eta19-phi3*/	3,1,2,2,1,3,7,13,5,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	5,11,0,1,11,1,1,11,2,3,27,1,4,27,2,1,
/* out0083_em-eta3-phi4*/	10,10,0,11,10,1,4,11,0,12,11,1,10,11,2,11,26,1,2,26,2,1,27,0,4,27,1,2,27,2,15,
/* out0084_em-eta4-phi4*/	4,9,1,13,10,0,5,10,2,5,26,2,13,
/* out0085_em-eta5-phi4*/	12,8,1,6,9,0,15,9,1,1,9,2,1,25,2,6,91,0,1,91,1,14,91,2,1,92,0,6,97,0,15,97,1,14,97,2,12,
/* out0086_em-eta6-phi4*/	9,8,0,12,8,1,9,8,2,4,82,0,9,82,1,7,91,1,2,91,2,5,92,0,2,92,2,3,
/* out0087_em-eta7-phi4*/	10,7,0,1,7,1,13,7,2,3,8,0,3,24,2,1,70,1,1,71,0,3,82,0,2,82,1,3,82,2,14,
/* out0088_em-eta8-phi4*/	6,6,1,2,7,0,10,7,2,5,70,1,5,71,0,10,71,2,4,
/* out0089_em-eta9-phi4*/	6,6,0,1,6,1,11,6,2,2,59,0,2,59,1,12,71,2,2,
/* out0090_em-eta10-phi4*/	6,4,5,4,6,2,10,66,0,1,48,0,2,59,1,4,59,2,7,
/* out0091_em-eta11-phi4*/	9,4,5,8,5,0,2,5,2,4,5,4,6,5,5,16,66,0,1,48,0,10,48,1,1,48,2,1,
/* out0092_em-eta12-phi4*/	8,4,3,1,5,2,8,5,3,13,5,4,8,47,0,1,47,1,1,36,1,1,48,2,8,
/* out0093_em-eta13-phi4*/	8,2,4,8,4,3,3,5,3,3,47,0,13,47,3,1,36,1,5,37,0,2,48,2,1,
/* out0094_em-eta14-phi4*/	8,2,4,2,2,5,15,3,5,1,47,3,4,36,1,2,36,2,1,37,0,2,37,2,1,
/* out0095_em-eta15-phi4*/	6,3,2,2,3,5,12,28,4,4,29,1,2,25,0,2,25,1,3,
/* out0096_em-eta16-phi4*/	5,3,2,1,28,1,5,29,1,10,25,0,1,25,1,3,
/* out0097_em-eta17-phi4*/	5,1,2,1,1,5,1,28,0,3,28,1,8,25,2,4,
/* out0098_em-eta18-phi4*/	4,1,2,6,13,2,1,28,0,4,25,2,2,
/* out0099_em-eta19-phi4*/	3,1,2,2,13,2,7,13,5,6,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	8,10,1,12,10,2,2,11,0,3,11,1,5,11,2,2,121,1,1,134,1,2,134,2,3,
/* out0104_em-eta4-phi5*/	5,9,1,2,9,2,5,10,2,9,121,0,10,121,1,11,
/* out0105_em-eta5-phi5*/	15,8,1,1,8,2,1,9,0,1,9,2,10,108,0,4,108,1,12,121,0,2,92,0,8,92,1,13,97,0,1,97,1,2,97,2,4,98,0,12,98,1,8,98,2,4,
/* out0106_em-eta6-phi5*/	8,8,2,10,95,0,4,95,1,4,108,0,8,82,1,3,83,0,9,92,1,3,92,2,13,
/* out0107_em-eta7-phi5*/	9,7,2,4,8,2,1,95,0,12,95,2,3,71,0,1,71,1,3,82,1,3,83,0,7,83,2,8,
/* out0108_em-eta8-phi5*/	7,7,2,4,83,0,9,83,1,4,95,2,1,71,0,2,71,1,13,71,2,5,
/* out0109_em-eta9-phi5*/	5,6,1,2,83,0,7,83,2,4,60,0,11,71,2,5,
/* out0110_em-eta10-phi5*/	6,6,2,1,66,0,7,66,1,3,48,1,1,60,0,5,60,2,7,
/* out0111_em-eta11-phi5*/	5,5,2,1,66,0,7,66,2,3,48,1,11,60,2,1,
/* out0112_em-eta12-phi5*/	8,5,2,3,47,1,11,48,0,2,48,1,12,66,2,1,37,0,1,48,1,3,48,2,5,
/* out0113_em-eta13-phi5*/	7,47,0,2,47,1,4,47,2,15,47,3,3,48,0,2,48,4,2,37,0,8,
/* out0114_em-eta14-phi5*/	6,47,2,1,47,3,8,48,3,12,48,4,2,37,0,3,37,2,4,
/* out0115_em-eta15-phi5*/	6,28,4,12,28,5,4,29,0,1,29,1,1,25,1,3,37,2,3,
/* out0116_em-eta16-phi5*/	4,28,2,4,29,0,11,29,1,2,25,1,5,
/* out0117_em-eta17-phi5*/	6,28,0,2,28,1,2,28,2,8,28,3,2,25,1,2,25,2,1,
/* out0118_em-eta18-phi5*/	4,13,2,2,28,0,7,28,3,2,25,2,1,
/* out0119_em-eta19-phi5*/	4,13,2,6,13,3,4,13,4,12,13,5,9,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	2,134,1,1,146,2,5,
/* out0123_em-eta3-phi6*/	7,121,1,1,134,1,13,134,2,13,135,0,10,135,1,4,146,1,4,146,2,8,
/* out0124_em-eta4-phi6*/	6,121,0,2,121,1,3,121,2,16,122,1,7,135,0,6,135,2,3,
/* out0125_em-eta5-phi6*/	14,108,1,4,108,2,12,109,1,2,121,0,2,122,0,8,122,1,2,93,0,13,93,1,8,98,0,4,98,1,8,98,2,12,99,0,4,99,1,2,99,2,1,
/* out0126_em-eta6-phi6*/	9,95,1,7,108,0,4,108,2,4,109,0,5,109,1,5,83,1,9,84,0,3,93,0,3,93,2,13,
/* out0127_em-eta7-phi6*/	9,95,1,5,95,2,11,96,1,4,109,0,1,72,0,3,72,1,1,83,1,7,83,2,8,84,0,3,
/* out0128_em-eta8-phi6*/	8,83,1,12,83,2,1,95,2,1,96,0,3,96,1,1,72,0,13,72,1,2,72,2,5,
/* out0129_em-eta9-phi6*/	5,66,1,1,83,2,11,84,0,3,60,1,11,72,2,5,
/* out0130_em-eta10-phi6*/	5,66,1,11,84,0,1,49,0,1,60,1,5,60,2,7,
/* out0131_em-eta11-phi6*/	4,66,2,10,67,0,1,49,0,11,60,2,1,
/* out0132_em-eta12-phi6*/	9,47,4,15,47,5,3,48,0,2,48,1,4,66,2,1,67,0,3,37,1,1,49,0,3,49,2,5,
/* out0133_em-eta13-phi6*/	5,47,5,5,48,0,10,48,4,9,48,5,4,37,1,8,
/* out0134_em-eta14-phi6*/	6,48,2,13,48,3,4,48,4,3,48,5,3,37,1,3,37,2,4,
/* out0135_em-eta15-phi6*/	5,28,5,12,29,0,1,29,5,6,26,0,3,37,2,3,
/* out0136_em-eta16-phi6*/	4,29,0,3,29,4,11,29,5,2,26,0,5,
/* out0137_em-eta17-phi6*/	6,28,2,4,28,3,2,29,3,3,29,4,5,26,0,2,26,2,1,
/* out0138_em-eta18-phi6*/	3,13,3,3,28,3,9,26,2,1,
/* out0139_em-eta19-phi6*/	5,12,0,12,12,2,16,12,3,5,13,3,8,13,4,4,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	4,146,1,3,146,2,3,147,0,1,147,1,4,
/* out0143_em-eta3-phi7*/	8,135,1,12,135,2,3,136,0,1,136,1,2,146,1,9,147,0,15,147,1,2,147,2,4,
/* out0144_em-eta4-phi7*/	4,122,1,6,122,2,7,135,2,10,136,0,13,
/* out0145_em-eta5-phi7*/	13,109,1,4,109,2,2,122,0,8,122,1,1,122,2,9,123,0,6,93,1,6,94,0,14,94,1,1,94,2,1,99,0,12,99,1,14,99,2,15,
/* out0146_em-eta6-phi7*/	9,109,0,7,109,1,5,109,2,13,84,0,7,84,1,9,93,1,2,93,2,3,94,0,2,94,2,5,
/* out0147_em-eta7-phi7*/	8,96,1,11,96,2,5,109,0,3,72,1,3,73,0,1,84,0,3,84,1,2,84,2,14,
/* out0148_em-eta8-phi7*/	6,84,1,2,96,0,13,96,2,2,72,1,10,72,2,4,73,0,5,
/* out0149_em-eta9-phi7*/	6,84,0,7,84,1,6,84,2,1,61,0,12,61,1,2,72,2,2,
/* out0150_em-eta10-phi7*/	7,66,1,1,68,1,4,84,0,5,84,2,5,49,1,2,61,0,4,61,2,7,
/* out0151_em-eta11-phi7*/	9,66,2,1,67,0,4,67,1,16,67,2,6,68,0,2,68,1,8,49,0,1,49,1,10,49,2,1,
/* out0152_em-eta12-phi7*/	8,47,4,1,47,5,2,67,0,8,67,2,8,67,3,13,68,3,1,38,0,1,49,2,8,
/* out0153_em-eta13-phi7*/	9,47,5,6,48,5,7,49,1,6,50,1,2,67,3,3,68,3,3,37,1,2,38,0,5,49,2,1,
/* out0154_em-eta14-phi7*/	9,48,2,3,48,5,2,49,0,9,49,1,9,49,2,1,37,1,2,37,2,1,38,0,2,38,2,1,
/* out0155_em-eta15-phi7*/	6,29,2,1,29,5,5,49,0,7,49,3,7,26,0,3,26,1,2,
/* out0156_em-eta16-phi7*/	6,29,2,11,29,3,1,29,5,3,49,3,1,26,0,3,26,1,1,
/* out0157_em-eta17-phi7*/	5,29,2,3,29,3,8,30,0,1,30,1,1,26,2,4,
/* out0158_em-eta18-phi7*/	6,12,3,1,13,3,1,28,3,1,29,3,4,30,0,6,26,2,2,
/* out0159_em-eta19-phi7*/	3,12,0,3,12,3,10,30,0,2,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	3,147,1,5,156,0,12,156,2,7,
/* out0163_em-eta3-phi8*/	6,136,1,6,147,1,5,147,2,12,148,0,7,148,1,12,156,0,3,
/* out0164_em-eta4-phi8*/	6,123,1,2,136,0,2,136,1,8,136,2,16,137,0,6,148,0,2,
/* out0165_em-eta5-phi8*/	8,123,0,8,123,1,13,123,2,9,94,1,15,94,2,2,95,0,13,95,1,2,95,2,1,
/* out0166_em-eta6-phi8*/	10,109,2,1,110,1,15,110,2,2,123,0,2,123,2,5,84,1,3,85,0,14,85,1,2,85,2,1,94,2,8,
/* out0167_em-eta7-phi8*/	10,96,2,5,97,1,2,110,0,13,110,1,1,73,0,5,73,1,7,84,1,2,84,2,2,85,0,2,85,2,5,
/* out0168_em-eta8-phi8*/	7,84,1,1,96,2,4,97,0,4,97,1,8,73,0,5,73,1,3,73,2,11,
/* out0169_em-eta9-phi8*/	7,84,1,7,84,2,4,85,1,1,97,0,3,61,1,13,62,0,2,73,2,2,
/* out0170_em-eta10-phi8*/	7,67,4,8,84,2,6,85,0,1,85,1,2,50,0,3,61,1,1,61,2,9,
/* out0171_em-eta11-phi8*/	9,67,2,1,67,4,8,67,5,9,68,0,14,68,1,4,68,4,2,68,5,1,49,1,3,50,0,8,
/* out0172_em-eta12-phi8*/	11,67,2,1,68,2,6,68,3,8,68,4,14,68,5,4,38,0,2,38,1,3,49,1,1,49,2,1,50,0,1,50,2,2,
/* out0173_em-eta13-phi8*/	7,49,4,6,50,0,1,50,1,14,68,2,3,68,3,4,38,0,5,38,1,2,
/* out0174_em-eta14-phi8*/	6,49,1,1,49,2,11,50,0,9,50,4,2,38,0,1,38,2,6,
/* out0175_em-eta15-phi8*/	6,49,2,4,49,3,6,50,3,5,50,4,4,26,1,4,38,2,1,
/* out0176_em-eta16-phi8*/	6,29,2,1,30,1,2,31,1,5,49,3,2,50,3,6,26,1,4,
/* out0177_em-eta17-phi8*/	4,30,1,11,30,2,1,31,1,2,26,2,4,
/* out0178_em-eta18-phi8*/	6,30,0,5,30,1,2,30,2,3,30,3,2,15,1,1,26,2,2,
/* out0179_em-eta19-phi8*/	3,12,0,1,30,0,2,30,3,7,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	5,156,0,1,156,2,9,157,0,10,157,1,12,157,2,3,
/* out0183_em-eta3-phi9*/	7,148,0,5,148,1,4,148,2,16,149,0,1,149,1,9,157,0,6,157,2,4,
/* out0184_em-eta4-phi9*/	5,137,0,7,137,1,16,137,2,9,148,0,2,149,0,3,
/* out0185_em-eta5-phi9*/	12,123,1,1,123,2,2,124,0,8,124,1,10,124,2,1,137,0,3,137,2,6,86,0,1,95,0,3,95,1,14,95,2,11,96,0,2,
/* out0186_em-eta6-phi9*/	9,110,2,9,111,0,1,111,1,2,124,0,8,124,2,4,85,1,14,85,2,2,86,0,9,95,2,4,
/* out0187_em-eta7-phi9*/	9,97,1,3,97,2,3,110,0,3,110,2,5,111,0,8,73,1,2,74,0,12,74,1,1,85,2,8,
/* out0188_em-eta8-phi9*/	9,97,0,3,97,1,3,97,2,11,62,0,3,62,1,3,73,1,4,73,2,3,74,0,3,74,2,3,
/* out0189_em-eta9-phi9*/	5,85,1,8,97,0,6,62,0,10,62,1,2,62,2,4,
/* out0190_em-eta10-phi9*/	7,85,0,6,85,1,5,85,2,1,50,0,2,50,1,7,62,0,1,62,2,4,
/* out0191_em-eta11-phi9*/	8,67,5,7,68,5,5,69,1,3,70,1,4,85,0,5,50,0,2,50,1,3,50,2,5,
/* out0192_em-eta12-phi9*/	7,68,2,6,68,5,6,69,0,9,69,1,12,38,1,3,39,0,1,50,2,6,
/* out0193_em-eta13-phi9*/	6,49,4,10,49,5,7,68,2,1,69,0,7,69,3,3,38,1,7,
/* out0194_em-eta14-phi9*/	6,49,5,6,50,0,6,50,4,6,50,5,5,27,0,1,38,2,6,
/* out0195_em-eta15-phi9*/	7,50,2,9,50,3,4,50,4,4,50,5,3,26,1,1,27,0,3,38,2,1,
/* out0196_em-eta16-phi9*/	6,30,4,6,31,1,6,50,2,2,50,3,1,26,1,3,27,0,2,
/* out0197_em-eta17-phi9*/	6,30,2,2,31,0,8,31,1,3,15,1,2,26,1,1,26,2,2,
/* out0198_em-eta18-phi9*/	5,30,2,8,30,3,3,31,0,1,31,4,2,15,1,4,
/* out0199_em-eta19-phi9*/	5,30,2,2,30,3,4,31,3,10,31,4,2,15,1,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	4,157,1,4,157,2,5,158,0,11,158,1,6,
/* out0203_em-eta3-phi10*/	7,149,0,3,149,1,7,149,2,15,150,1,4,157,2,4,158,0,5,158,2,12,
/* out0204_em-eta4-phi10*/	8,137,2,1,138,0,1,138,1,15,138,2,7,149,0,9,149,2,1,150,0,1,150,1,1,
/* out0205_em-eta5-phi10*/	11,124,1,6,124,2,4,125,0,3,125,1,3,138,0,13,138,1,1,86,0,1,86,1,7,87,0,1,96,0,14,96,2,14,
/* out0206_em-eta6-phi10*/	7,111,1,11,124,2,7,125,0,8,75,0,1,86,0,5,86,1,8,86,2,14,
/* out0207_em-eta7-phi10*/	8,111,0,6,111,1,3,111,2,12,74,0,1,74,1,15,74,2,3,75,0,3,86,2,1,
/* out0208_em-eta8-phi10*/	7,97,2,2,98,1,13,111,0,1,111,2,1,62,1,4,63,0,6,74,2,10,
/* out0209_em-eta9-phi10*/	7,85,2,6,98,0,7,98,1,1,51,0,1,62,1,7,62,2,5,63,0,2,
/* out0210_em-eta10-phi10*/	6,85,0,1,85,2,9,86,1,1,50,1,2,51,0,9,62,2,3,
/* out0211_em-eta11-phi10*/	11,69,4,12,69,5,1,70,0,2,70,1,11,85,0,3,39,0,1,39,1,1,50,1,4,50,2,2,51,0,3,51,2,1,
/* out0212_em-eta12-phi10*/	7,69,1,1,69,2,14,70,0,11,70,1,1,70,4,6,39,0,8,50,2,1,
/* out0213_em-eta13-phi10*/	8,49,5,1,69,2,2,69,3,13,70,3,9,70,4,2,38,1,1,39,0,5,39,2,2,
/* out0214_em-eta14-phi10*/	8,49,5,2,50,5,7,51,1,9,52,1,4,70,3,1,27,0,3,27,1,3,38,2,1,
/* out0215_em-eta15-phi10*/	5,50,2,5,50,5,1,51,0,10,51,1,3,27,0,5,
/* out0216_em-eta16-phi10*/	5,30,4,10,30,5,2,51,0,4,27,0,2,27,2,2,
/* out0217_em-eta17-phi10*/	5,30,5,6,31,0,7,31,4,1,15,2,3,27,2,2,
/* out0218_em-eta18-phi10*/	5,31,2,1,31,4,10,31,5,1,15,1,3,15,2,2,
/* out0219_em-eta19-phi10*/	4,31,2,2,31,3,6,31,4,1,15,1,2,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	1,158,1,6,
/* out0223_em-eta3-phi11*/	8,150,0,1,150,1,11,150,2,14,158,1,4,158,2,4,159,0,12,159,1,8,159,2,4,
/* out0224_em-eta4-phi11*/	4,138,2,7,139,1,13,150,0,14,150,2,2,
/* out0225_em-eta5-phi11*/	10,125,1,13,125,2,3,138,0,2,138,2,2,139,0,8,139,1,3,87,0,11,87,1,12,87,2,3,96,2,2,
/* out0226_em-eta6-phi11*/	9,112,1,5,125,0,5,125,2,13,75,0,4,75,1,10,86,1,1,86,2,1,87,0,4,87,2,9,
/* out0227_em-eta7-phi11*/	9,98,1,1,98,2,1,111,2,3,112,0,14,112,1,3,63,1,1,75,0,8,75,1,2,75,2,12,
/* out0228_em-eta8-phi11*/	7,98,0,1,98,1,1,98,2,13,112,0,2,63,0,6,63,1,11,63,2,3,
/* out0229_em-eta9-phi11*/	6,86,1,5,98,0,8,98,2,2,51,1,5,63,0,2,63,2,9,
/* out0230_em-eta10-phi11*/	5,86,0,2,86,1,10,51,0,3,51,1,7,51,2,3,
/* out0231_em-eta11-phi11*/	5,69,4,4,69,5,12,86,0,6,39,1,3,51,2,8,
/* out0232_em-eta12-phi11*/	8,69,5,3,70,0,3,70,2,4,70,4,7,70,5,16,39,0,1,39,1,8,39,2,1,
/* out0233_em-eta13-phi11*/	6,51,4,7,52,1,2,70,2,12,70,3,6,70,4,1,39,2,8,
/* out0234_em-eta14-phi11*/	7,51,1,2,51,2,2,51,4,1,52,0,8,52,1,10,27,1,5,39,2,1,
/* out0235_em-eta15-phi11*/	6,51,0,1,51,1,2,51,2,14,51,3,2,27,1,4,27,2,2,
/* out0236_em-eta16-phi11*/	4,30,5,2,51,0,1,51,3,13,27,2,5,
/* out0237_em-eta17-phi11*/	5,30,5,6,31,5,7,51,3,1,15,2,3,27,2,2,
/* out0238_em-eta18-phi11*/	3,31,2,4,31,5,8,15,2,4,
/* out0239_em-eta19-phi11*/	2,31,2,9,15,1,2,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	2,160,0,8,160,1,3,
/* out0243_em-eta3-phi12*/	8,151,0,6,151,1,15,151,2,4,159,0,4,159,1,8,159,2,12,160,0,8,160,2,5,
/* out0244_em-eta4-phi12*/	4,139,2,13,140,1,7,151,0,10,151,2,7,
/* out0245_em-eta5-phi12*/	12,126,1,10,126,2,5,139,0,8,139,2,3,140,0,2,140,1,2,76,0,1,76,1,4,87,1,4,87,2,2,88,0,15,88,2,8,
/* out0246_em-eta6-phi12*/	9,112,1,5,126,0,12,126,1,6,126,2,1,75,1,2,76,0,15,76,1,4,76,2,5,87,2,2,
/* out0247_em-eta7-phi12*/	9,99,1,1,112,1,3,112,2,14,113,0,3,64,0,9,64,1,6,75,1,2,75,2,4,76,2,2,
/* out0248_em-eta8-phi12*/	9,99,0,6,99,1,9,112,2,2,52,0,1,52,1,2,63,1,4,63,2,2,64,0,7,64,2,4,
/* out0249_em-eta9-phi12*/	6,86,2,5,99,0,10,51,1,1,52,0,12,52,1,1,63,2,2,
/* out0250_em-eta10-phi12*/	8,86,0,2,86,2,10,40,0,1,40,1,2,51,1,3,51,2,2,52,0,3,52,2,2,
/* out0251_em-eta11-phi12*/	5,71,4,7,71,5,9,86,0,6,40,0,9,51,2,2,
/* out0252_em-eta12-phi12*/	10,71,2,1,71,4,9,71,5,1,72,0,9,72,1,12,28,1,1,39,1,4,39,2,1,40,0,4,40,2,1,
/* out0253_em-eta13-phi12*/	7,51,4,7,51,5,2,71,0,1,71,1,13,72,1,4,28,0,5,39,2,3,
/* out0254_em-eta14-phi12*/	7,51,4,1,51,5,10,52,0,8,52,4,2,52,5,2,27,1,1,28,0,5,
/* out0255_em-eta15-phi12*/	7,52,2,1,52,3,2,52,4,14,52,5,2,27,1,3,27,2,1,28,0,1,
/* out0256_em-eta16-phi12*/	5,32,4,2,52,2,1,52,3,13,16,0,2,27,2,2,
/* out0257_em-eta17-phi12*/	3,32,4,12,52,3,1,16,0,3,
/* out0258_em-eta18-phi12*/	4,32,4,2,33,1,10,15,2,3,16,0,1,
/* out0259_em-eta19-phi12*/	4,32,1,5,33,1,5,15,1,1,15,2,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	3,160,1,10,161,0,6,161,1,5,
/* out0263_em-eta3-phi13*/	8,151,1,1,151,2,3,152,0,8,152,1,14,152,2,2,160,1,3,160,2,11,161,0,5,
/* out0264_em-eta4-phi13*/	7,140,0,1,140,1,7,140,2,15,141,0,1,151,2,2,152,0,8,152,2,2,
/* out0265_em-eta5-phi13*/	10,126,2,6,127,1,10,140,0,13,140,2,1,76,1,2,77,0,14,77,1,7,77,2,1,88,0,1,88,2,8,
/* out0266_em-eta6-phi13*/	11,113,1,11,126,0,4,126,2,4,127,0,3,127,1,3,65,0,6,65,1,2,76,1,6,76,2,8,77,0,2,77,2,3,
/* out0267_em-eta7-phi13*/	8,113,0,12,113,1,3,113,2,6,64,1,10,64,2,3,65,0,8,65,2,1,76,2,1,
/* out0268_em-eta8-phi13*/	9,99,1,6,99,2,8,100,0,2,100,1,1,113,0,1,113,2,1,52,1,4,53,0,7,64,2,9,
/* out0269_em-eta9-phi13*/	4,87,1,6,99,2,8,52,1,9,52,2,7,
/* out0270_em-eta10-phi13*/	6,86,2,1,87,0,1,87,1,9,40,1,6,41,0,1,52,2,6,
/* out0271_em-eta11-phi13*/	9,71,5,6,72,0,1,72,2,3,72,4,1,72,5,16,87,0,3,40,0,2,40,1,6,40,2,3,
/* out0272_em-eta12-phi13*/	6,71,2,10,72,0,6,72,3,1,72,4,15,28,1,2,40,2,7,
/* out0273_em-eta13-phi13*/	7,53,4,1,71,0,14,71,1,3,71,2,5,71,3,5,28,0,2,28,1,6,
/* out0274_em-eta14-phi13*/	7,51,5,4,52,5,9,53,4,9,54,1,1,71,0,1,28,0,3,28,2,3,
/* out0275_em-eta15-phi13*/	5,52,2,10,52,5,3,54,1,5,16,1,2,28,2,3,
/* out0276_em-eta16-phi13*/	5,32,5,10,33,5,2,52,2,4,16,0,3,16,1,2,
/* out0277_em-eta17-phi13*/	3,32,5,6,33,0,7,16,0,4,
/* out0278_em-eta18-phi13*/	5,32,2,3,33,0,7,33,1,1,16,0,2,16,2,1,
/* out0279_em-eta19-phi13*/	5,32,0,10,32,1,8,32,2,2,16,0,1,16,2,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	5,161,0,1,161,1,11,161,2,11,162,0,9,162,2,1,
/* out0283_em-eta3-phi14*/	6,152,1,2,152,2,8,153,0,13,153,1,12,161,0,4,161,2,5,
/* out0284_em-eta4-phi14*/	5,141,0,9,141,1,16,141,2,7,152,2,4,153,0,2,
/* out0285_em-eta5-phi14*/	13,127,0,1,127,1,3,127,2,15,128,1,3,141,0,6,141,2,3,66,0,5,66,1,2,77,1,9,77,2,8,78,0,14,78,1,13,78,2,12,
/* out0286_em-eta6-phi14*/	10,113,1,2,113,2,1,114,1,9,127,0,12,127,2,1,65,0,1,65,1,14,65,2,2,66,0,8,77,2,4,
/* out0287_em-eta7-phi14*/	8,100,1,5,113,2,8,114,0,3,114,1,5,53,1,7,54,0,2,65,0,1,65,2,13,
/* out0288_em-eta8-phi14*/	6,100,0,8,100,1,7,100,2,2,53,0,7,53,1,7,53,2,6,
/* out0289_em-eta9-phi14*/	7,87,2,8,100,0,6,41,0,3,41,1,6,52,2,1,53,0,2,53,2,4,
/* out0290_em-eta10-phi14*/	6,87,0,6,87,1,1,87,2,5,41,0,11,41,1,1,41,2,2,
/* out0291_em-eta11-phi14*/	9,72,2,8,73,4,12,87,0,5,29,0,2,29,1,1,40,1,2,40,2,3,41,0,1,41,2,1,
/* out0292_em-eta12-phi14*/	8,71,3,2,72,2,5,72,3,15,73,4,3,74,1,9,28,1,1,29,0,7,40,2,2,
/* out0293_em-eta13-phi14*/	8,53,4,2,53,5,13,54,5,2,71,3,9,73,1,1,28,1,6,28,2,1,29,0,1,
/* out0294_em-eta14-phi14*/	5,53,4,4,53,5,3,54,0,12,54,1,4,28,2,6,
/* out0295_em-eta15-phi14*/	7,53,1,9,53,2,2,54,0,2,54,1,6,16,1,3,17,0,1,28,2,2,
/* out0296_em-eta16-phi14*/	4,33,2,1,33,5,11,53,1,4,16,1,5,
/* out0297_em-eta17-phi14*/	5,33,0,1,33,4,10,33,5,3,16,1,1,16,2,3,
/* out0298_em-eta18-phi14*/	4,32,2,7,33,0,1,33,4,3,16,2,3,
/* out0299_em-eta19-phi14*/	5,32,0,4,32,1,3,32,2,3,32,3,2,16,2,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	4,154,1,3,154,2,2,162,0,5,162,2,14,
/* out0303_em-eta3-phi15*/	7,142,1,6,153,1,4,153,2,15,154,0,4,154,1,13,162,0,2,162,2,1,
/* out0304_em-eta4-phi15*/	8,128,1,1,128,2,2,141,2,6,142,0,16,142,1,8,142,2,2,153,0,1,153,2,1,
/* out0305_em-eta5-phi15*/	11,128,0,8,128,1,12,128,2,10,66,1,14,66,2,2,67,0,16,67,1,10,67,2,1,78,0,2,78,1,3,78,2,4,
/* out0306_em-eta6-phi15*/	9,114,1,2,114,2,15,115,1,1,128,0,6,54,0,1,54,1,8,55,0,2,66,0,3,66,2,14,
/* out0307_em-eta7-phi15*/	7,100,1,2,101,1,4,114,0,13,114,2,1,54,0,12,54,1,5,54,2,6,
/* out0308_em-eta8-phi15*/	11,88,1,1,88,2,1,100,1,1,100,2,11,101,1,4,42,0,6,42,1,4,53,1,2,53,2,5,54,0,1,54,2,2,
/* out0309_em-eta9-phi15*/	6,87,2,1,88,1,10,100,2,3,41,1,8,42,0,7,53,2,1,
/* out0310_em-eta10-phi15*/	9,73,5,3,74,5,5,87,0,1,87,2,2,88,0,3,88,1,4,30,0,1,41,1,1,41,2,11,
/* out0311_em-eta11-phi15*/	8,73,4,1,73,5,13,74,0,10,74,1,1,74,4,7,74,5,7,29,1,9,41,2,2,
/* out0312_em-eta12-phi15*/	8,73,0,1,73,1,11,73,2,9,74,0,6,74,1,6,29,0,4,29,1,2,29,2,4,
/* out0313_em-eta13-phi15*/	8,54,2,6,54,4,1,54,5,14,73,0,3,73,1,4,17,1,2,29,0,2,29,2,3,
/* out0314_em-eta14-phi15*/	7,53,2,5,54,0,2,54,3,1,54,4,15,17,0,5,17,1,1,28,2,1,
/* out0315_em-eta15-phi15*/	5,53,0,5,53,1,3,53,2,9,53,3,3,17,0,5,
/* out0316_em-eta16-phi15*/	6,33,2,7,34,1,1,35,1,1,53,0,8,16,1,3,17,0,1,
/* out0317_em-eta17-phi15*/	4,33,2,7,33,3,6,33,4,1,16,2,4,
/* out0318_em-eta18-phi15*/	5,32,2,1,32,3,3,33,3,5,33,4,2,16,2,3,
/* out0319_em-eta19-phi15*/	3,14,4,1,32,0,2,32,3,7,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	4,154,2,6,155,0,1,155,1,1,155,2,3,
/* out0323_em-eta3-phi16*/	9,142,1,2,142,2,1,143,1,11,143,2,4,154,0,12,154,2,8,155,0,12,155,1,10,155,2,11,
/* out0324_em-eta4-phi16*/	5,129,1,7,129,2,6,142,2,13,143,0,5,143,1,5,
/* out0325_em-eta5-phi16*/	13,115,1,2,115,2,4,128,0,2,128,2,4,129,0,8,129,1,9,129,2,1,55,0,1,55,1,10,56,0,5,56,1,6,67,1,6,67,2,15,
/* out0326_em-eta6-phi16*/	8,115,0,7,115,1,13,115,2,5,43,1,1,54,1,1,55,0,13,55,1,4,55,2,10,
/* out0327_em-eta7-phi16*/	7,101,1,5,101,2,11,115,0,3,43,0,10,43,1,3,54,1,2,54,2,8,
/* out0328_em-eta8-phi16*/	7,88,2,2,101,0,13,101,1,3,42,0,1,42,1,12,42,2,4,43,0,2,
/* out0329_em-eta9-phi16*/	6,88,0,2,88,1,1,88,2,11,30,1,4,42,0,2,42,2,10,
/* out0330_em-eta10-phi16*/	6,74,2,3,74,5,1,75,1,1,88,0,10,30,0,9,30,1,4,
/* out0331_em-eta11-phi16*/	8,74,2,13,74,3,12,74,4,8,74,5,3,75,1,1,29,1,4,30,0,6,30,2,1,
/* out0332_em-eta12-phi16*/	9,55,4,1,56,1,2,73,0,6,73,2,7,73,3,14,74,3,2,74,4,1,18,0,2,29,2,7,
/* out0333_em-eta13-phi16*/	7,54,2,8,55,1,7,56,1,6,73,0,6,17,1,5,18,0,1,29,2,2,
/* out0334_em-eta14-phi16*/	8,53,3,1,54,2,2,54,3,15,55,0,3,55,1,2,17,0,1,17,1,4,17,2,1,
/* out0335_em-eta15-phi16*/	6,34,4,4,35,1,2,53,0,2,53,3,12,17,0,2,17,2,3,
/* out0336_em-eta16-phi16*/	6,34,1,5,35,1,10,53,0,1,7,2,1,17,0,1,17,2,2,
/* out0337_em-eta17-phi16*/	5,33,2,1,33,3,1,34,0,3,34,1,8,7,1,3,
/* out0338_em-eta18-phi16*/	6,14,5,1,15,5,1,32,3,2,33,3,4,34,0,4,7,1,3,
/* out0339_em-eta19-phi16*/	3,14,4,3,14,5,10,32,3,2,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	8,130,1,1,143,0,2,143,2,12,144,0,3,144,2,2,155,0,3,155,1,5,155,2,2,
/* out0344_em-eta4-phi17*/	4,129,2,7,130,0,10,130,1,11,143,0,9,
/* out0345_em-eta5-phi17*/	11,115,2,2,116,0,4,116,1,12,129,0,8,129,2,2,130,0,2,44,1,5,55,1,1,56,0,11,56,1,10,56,2,16,
/* out0346_em-eta6-phi17*/	9,102,1,7,115,0,5,115,2,5,116,0,8,43,1,3,44,0,15,44,1,3,55,1,1,55,2,6,
/* out0347_em-eta7-phi17*/	8,101,2,4,102,0,11,102,1,5,115,0,1,43,0,2,43,1,9,43,2,11,44,0,1,
/* out0348_em-eta8-phi17*/	10,89,1,9,89,2,4,101,0,3,101,2,1,102,0,1,31,0,4,31,1,8,42,2,1,43,0,2,43,2,5,
/* out0349_em-eta9-phi17*/	6,88,2,2,89,0,4,89,1,7,30,1,3,31,0,12,42,2,1,
/* out0350_em-eta10-phi17*/	5,75,1,7,75,2,3,88,0,1,30,1,5,30,2,9,
/* out0351_em-eta11-phi17*/	5,74,3,1,75,0,3,75,1,7,18,1,5,30,2,6,
/* out0352_em-eta12-phi17*/	9,55,4,15,55,5,4,56,0,2,56,1,3,73,3,2,74,3,1,75,0,1,18,0,7,18,1,3,
/* out0353_em-eta13-phi17*/	6,55,1,4,55,2,9,56,0,10,56,1,5,17,1,2,18,0,6,
/* out0354_em-eta14-phi17*/	6,55,0,13,55,1,3,55,2,3,55,3,4,17,1,2,17,2,4,
/* out0355_em-eta15-phi17*/	5,34,4,12,34,5,4,35,0,1,35,1,1,17,2,5,
/* out0356_em-eta16-phi17*/	5,34,2,4,35,0,11,35,1,2,7,2,4,17,2,1,
/* out0357_em-eta17-phi17*/	6,34,0,2,34,1,2,34,2,8,34,3,2,7,1,2,7,2,2,
/* out0358_em-eta18-phi17*/	4,15,5,3,34,0,7,34,3,2,7,1,3,
/* out0359_em-eta19-phi17*/	5,14,4,12,14,5,5,15,0,16,15,4,4,15,5,8,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	3,144,2,1,145,0,1,145,2,4,
/* out0363_em-eta3-phi18*/	6,130,1,1,131,1,10,131,2,4,144,0,13,144,2,13,145,0,12,
/* out0364_em-eta4-phi18*/	7,117,1,5,117,2,2,130,0,2,130,1,3,130,2,16,131,0,3,131,1,6,
/* out0365_em-eta5-phi18*/	12,103,1,1,103,2,1,116,1,4,116,2,12,117,0,1,117,1,10,130,0,2,33,1,1,44,1,5,45,0,16,45,1,15,45,2,9,
/* out0366_em-eta6-phi18*/	10,102,1,4,102,2,4,103,1,10,116,0,4,116,2,4,32,1,3,33,0,6,33,1,1,44,1,3,44,2,15,
/* out0367_em-eta7-phi18*/	8,90,1,4,102,0,3,102,2,12,103,1,1,32,0,11,32,1,9,32,2,2,44,2,1,
/* out0368_em-eta8-phi18*/	9,89,0,1,89,2,12,90,1,4,102,0,1,20,0,1,31,1,8,31,2,4,32,0,5,32,2,2,
/* out0369_em-eta9-phi18*/	6,75,2,1,76,1,3,89,0,11,19,1,3,20,0,1,31,2,12,
/* out0370_em-eta10-phi18*/	4,75,2,11,76,1,1,19,0,9,19,1,5,
/* out0371_em-eta11-phi18*/	4,57,4,1,75,0,10,18,1,5,19,0,6,
/* out0372_em-eta12-phi18*/	7,55,5,12,56,0,2,56,5,11,57,4,3,75,0,1,18,1,3,18,2,7,
/* out0373_em-eta13-phi18*/	8,55,2,2,56,0,2,56,2,2,56,3,3,56,4,15,56,5,4,8,1,2,18,2,6,
/* out0374_em-eta14-phi18*/	6,55,2,2,55,3,12,56,3,8,56,4,1,8,0,4,8,1,2,
/* out0375_em-eta15-phi18*/	4,34,5,12,35,0,1,35,5,6,8,0,5,
/* out0376_em-eta16-phi18*/	5,35,0,3,35,4,11,35,5,2,7,2,4,8,0,1,
/* out0377_em-eta17-phi18*/	7,34,2,4,34,3,2,35,3,3,35,4,5,7,0,2,7,1,1,7,2,3,
/* out0378_em-eta18-phi18*/	3,15,2,2,34,3,9,7,1,3,
/* out0379_em-eta19-phi18*/	4,15,2,6,15,3,9,15,4,12,15,5,4,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	2,132,1,6,145,2,6,
/* out0383_em-eta3-phi19*/	8,118,1,1,118,2,2,131,0,3,131,2,12,132,0,12,132,1,8,145,0,3,145,2,6,
/* out0384_em-eta4-phi19*/	3,117,2,13,118,1,13,131,0,10,
/* out0385_em-eta5-phi19*/	13,103,2,6,104,0,2,104,1,4,117,0,15,117,1,1,117,2,1,33,1,10,33,2,1,34,0,16,34,1,12,34,2,2,45,1,1,45,2,7,
/* out0386_em-eta6-phi19*/	8,103,0,12,103,1,4,103,2,9,21,1,1,32,1,1,33,0,10,33,1,4,33,2,13,
/* out0387_em-eta7-phi19*/	8,90,0,1,90,1,3,90,2,13,103,0,3,21,0,8,21,1,2,32,1,3,32,2,10,
/* out0388_em-eta8-phi19*/	7,76,2,2,90,0,10,90,1,5,20,0,4,20,1,12,20,2,1,32,2,2,
/* out0389_em-eta9-phi19*/	6,76,0,1,76,1,7,76,2,6,19,1,4,20,0,10,20,2,2,
/* out0390_em-eta10-phi19*/	6,58,5,4,75,2,1,76,0,5,76,1,5,19,1,4,19,2,9,
/* out0391_em-eta11-phi19*/	9,57,4,4,57,5,16,58,0,6,58,4,2,58,5,8,75,0,1,9,1,4,19,0,1,19,2,6,
/* out0392_em-eta12-phi19*/	8,56,2,1,56,5,1,57,1,1,57,4,8,58,0,8,58,1,13,9,0,7,18,2,2,
/* out0393_em-eta13-phi19*/	9,36,5,6,37,5,2,56,2,13,56,3,1,57,1,3,58,1,3,8,1,5,9,0,2,18,2,1,
/* out0394_em-eta14-phi19*/	7,36,4,9,36,5,9,37,0,1,56,3,4,8,0,1,8,1,4,8,2,1,
/* out0395_em-eta15-phi19*/	6,35,2,1,35,5,5,36,4,7,37,1,7,8,0,3,8,2,2,
/* out0396_em-eta16-phi19*/	8,35,2,11,35,3,1,35,5,3,37,1,1,7,0,1,7,2,2,8,0,2,8,2,1,
/* out0397_em-eta17-phi19*/	5,16,4,1,16,5,1,35,2,3,35,3,8,7,0,8,
/* out0398_em-eta18-phi19*/	6,15,2,1,16,4,6,34,3,1,35,3,4,7,0,4,7,1,1,
/* out0399_em-eta19-phi19*/	3,15,2,7,15,3,6,16,4,2,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	4,132,1,2,132,2,3,133,0,14,133,2,5,
/* out0403_em-eta3-phi20*/	7,118,2,6,119,1,15,119,2,4,132,0,4,132,2,13,133,0,1,133,2,2,
/* out0404_em-eta4-phi20*/	8,104,1,2,104,2,1,105,1,6,118,0,16,118,1,2,118,2,8,119,0,1,119,1,1,
/* out0405_em-eta5-phi20*/	10,104,0,8,104,1,10,104,2,12,22,0,2,22,1,14,23,0,4,23,1,3,23,2,2,34,1,4,34,2,14,
/* out0406_em-eta6-phi20*/	9,91,1,15,91,2,2,103,0,1,104,0,6,21,1,8,21,2,1,22,0,14,22,2,3,33,2,2,
/* out0407_em-eta7-phi20*/	8,77,2,2,90,0,1,90,2,3,91,0,13,91,1,1,21,0,6,21,1,5,21,2,12,
/* out0408_em-eta8-phi20*/	10,76,2,1,77,1,11,77,2,1,90,0,4,11,0,5,11,1,2,20,1,4,20,2,6,21,0,2,21,2,1,
/* out0409_em-eta9-phi20*/	7,59,1,1,76,0,4,76,2,7,77,1,3,10,1,8,11,0,1,20,2,7,
/* out0410_em-eta10-phi20*/	7,58,2,8,59,0,1,59,1,2,76,0,6,10,0,11,10,1,1,19,2,1,
/* out0411_em-eta11-phi20*/	9,57,2,2,57,3,1,58,0,1,58,2,8,58,3,9,58,4,14,58,5,4,9,1,9,10,0,2,
/* out0412_em-eta12-phi20*/	8,57,0,6,57,1,8,57,2,14,57,3,4,58,0,1,9,0,4,9,1,2,9,2,4,
/* out0413_em-eta13-phi20*/	8,37,2,6,37,4,1,37,5,14,57,0,3,57,1,4,8,1,2,9,0,3,9,2,2,
/* out0414_em-eta14-phi20*/	7,36,2,2,36,5,1,37,0,11,37,4,9,1,0,1,8,1,1,8,2,5,
/* out0415_em-eta15-phi20*/	5,36,1,5,36,2,4,37,0,4,37,1,6,8,2,5,
/* out0416_em-eta16-phi20*/	7,16,5,2,17,5,5,35,2,1,36,1,6,37,1,2,0,1,3,8,2,1,
/* out0417_em-eta17-phi20*/	4,16,5,11,17,0,1,17,5,2,0,0,4,
/* out0418_em-eta18-phi20*/	6,16,4,5,16,5,2,17,0,3,17,1,2,0,0,3,7,0,1,
/* out0419_em-eta19-phi20*/	3,15,3,1,16,4,2,17,1,7,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	5,120,0,16,120,1,8,120,2,3,133,0,1,133,2,9,
/* out0423_em-eta3-phi21*/	5,106,1,8,106,2,2,119,0,13,119,2,12,120,2,11,
/* out0424_em-eta4-phi21*/	5,105,0,9,105,1,7,105,2,16,106,1,4,119,0,2,
/* out0425_em-eta5-phi21*/	13,92,0,1,92,1,15,92,2,3,104,2,3,105,0,6,105,1,3,13,0,8,13,1,9,22,1,2,22,2,5,23,0,12,23,1,13,23,2,14,
/* out0426_em-eta6-phi21*/	10,78,1,1,78,2,2,91,2,9,92,0,12,92,1,1,12,0,2,12,1,14,12,2,1,13,0,4,22,2,8,
/* out0427_em-eta7-phi21*/	8,77,2,5,78,1,8,91,0,3,91,2,5,11,1,7,12,0,13,12,2,1,21,2,2,
/* out0428_em-eta8-phi21*/	6,77,0,8,77,1,2,77,2,7,11,0,6,11,1,7,11,2,7,
/* out0429_em-eta9-phi21*/	7,59,1,8,77,0,6,3,0,1,10,1,6,10,2,3,11,0,4,11,2,2,
/* out0430_em-eta10-phi21*/	6,59,0,6,59,1,5,59,2,1,10,0,2,10,1,1,10,2,11,
/* out0431_em-eta11-phi21*/	10,38,4,8,57,3,5,58,3,7,59,0,5,2,0,3,2,1,2,9,1,1,9,2,2,10,0,1,10,2,1,
/* out0432_em-eta12-phi21*/	8,38,1,2,38,4,5,39,1,15,57,0,6,57,3,6,1,1,1,2,0,2,9,2,7,
/* out0433_em-eta13-phi21*/	7,37,2,10,37,3,7,38,1,9,57,0,1,1,0,1,1,1,6,9,2,1,
/* out0434_em-eta14-phi21*/	5,36,2,6,36,3,5,37,3,6,37,4,6,1,0,6,
/* out0435_em-eta15-phi21*/	7,36,0,9,36,1,4,36,2,4,36,3,3,0,1,3,1,0,2,8,2,1,
/* out0436_em-eta16-phi21*/	5,17,2,6,17,5,6,36,0,2,36,1,1,0,1,5,
/* out0437_em-eta17-phi21*/	5,17,0,2,17,4,8,17,5,3,0,0,3,0,1,1,
/* out0438_em-eta18-phi21*/	5,16,2,2,17,0,8,17,1,3,17,4,1,0,0,3,
/* out0439_em-eta19-phi21*/	5,16,1,10,16,2,2,17,0,2,17,1,4,0,0,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	3,107,0,5,107,1,11,120,1,7,
/* out0443_em-eta3-phi22*/	9,94,1,3,94,2,1,106,0,8,106,1,2,106,2,14,107,0,11,107,2,4,120,1,1,120,2,2,
/* out0444_em-eta4-phi22*/	7,93,0,1,93,1,15,93,2,7,94,1,2,105,0,1,106,0,8,106,1,2,
/* out0445_em-eta5-phi22*/	10,79,1,6,92,2,10,93,0,13,93,1,1,5,1,2,6,0,8,6,2,1,13,0,1,13,1,7,13,2,14,
/* out0446_em-eta6-phi22*/	11,78,2,11,79,0,4,79,1,4,92,0,3,92,2,3,5,0,8,5,1,6,12,1,2,12,2,6,13,0,3,13,2,2,
/* out0447_em-eta7-phi22*/	8,78,0,12,78,1,6,78,2,3,4,0,3,4,1,10,5,0,1,12,0,1,12,2,8,
/* out0448_em-eta8-phi22*/	9,60,1,8,60,2,6,77,0,2,77,2,1,78,0,1,78,1,1,3,1,4,4,0,9,11,2,7,
/* out0449_em-eta9-phi22*/	4,59,2,6,60,1,8,3,0,7,3,1,9,
/* out0450_em-eta10-phi22*/	6,40,1,1,59,0,1,59,2,9,2,1,6,3,0,6,10,2,1,
/* out0451_em-eta11-phi22*/	10,38,4,3,38,5,16,39,0,1,39,4,1,39,5,6,40,0,8,59,0,3,2,0,3,2,1,6,2,2,2,
/* out0452_em-eta12-phi22*/	6,38,2,10,39,0,15,39,1,1,39,4,6,1,1,2,2,0,7,
/* out0453_em-eta13-phi22*/	7,37,3,1,38,0,14,38,1,5,38,2,5,38,3,3,1,1,6,1,2,2,
/* out0454_em-eta14-phi22*/	7,18,5,9,19,5,4,36,3,7,37,3,2,38,0,1,1,0,3,1,2,3,
/* out0455_em-eta15-phi22*/	6,18,4,10,18,5,3,36,0,5,36,3,1,0,1,2,1,0,3,
/* out0456_em-eta16-phi22*/	5,17,2,10,17,3,2,18,4,4,0,1,2,0,2,3,
/* out0457_em-eta17-phi22*/	4,16,2,1,17,3,6,17,4,7,0,2,4,
/* out0458_em-eta18-phi22*/	5,16,0,1,16,2,10,16,3,1,0,0,1,0,2,2,
/* out0459_em-eta19-phi22*/	5,16,0,2,16,1,6,16,2,1,0,0,1,0,2,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	2,107,1,5,107,2,4,
/* out0463_em-eta3-phi23*/	4,94,0,6,94,1,4,94,2,15,107,2,8,
/* out0464_em-eta4-phi23*/	5,80,0,8,80,1,13,93,2,7,94,0,10,94,1,7,
/* out0465_em-eta5-phi23*/	10,79,1,5,79,2,10,80,0,8,80,1,3,93,0,2,93,2,2,5,1,4,5,2,1,6,0,8,6,2,15,
/* out0466_em-eta6-phi23*/	7,61,2,13,79,0,12,79,1,1,79,2,6,5,0,5,5,1,4,5,2,15,
/* out0467_em-eta7-phi23*/	7,60,2,1,61,1,14,61,2,3,78,0,3,4,1,6,4,2,9,5,0,2,
/* out0468_em-eta8-phi23*/	7,60,0,6,60,2,9,61,1,2,3,1,2,3,2,1,4,0,4,4,2,7,
/* out0469_em-eta9-phi23*/	5,40,1,5,40,2,1,60,0,10,3,1,1,3,2,12,
/* out0470_em-eta10-phi23*/	7,40,0,2,40,1,10,40,2,15,2,1,2,2,2,1,3,0,2,3,2,3,
/* out0471_em-eta11-phi23*/	4,39,2,7,39,5,9,40,0,6,2,2,9,
/* out0472_em-eta12-phi23*/	8,38,2,1,39,2,9,39,3,12,39,4,9,39,5,1,1,1,1,2,0,1,2,2,4,
/* out0473_em-eta13-phi23*/	6,19,2,7,19,5,2,38,0,1,38,3,13,39,3,4,1,2,5,
/* out0474_em-eta14-phi23*/	6,18,5,2,19,0,2,19,2,9,19,4,8,19,5,10,1,2,5,
/* out0475_em-eta15-phi23*/	6,18,4,1,18,5,2,19,0,14,19,1,2,19,4,8,1,2,1,
/* out0476_em-eta16-phi23*/	4,17,3,2,18,4,1,19,1,13,0,2,2,
/* out0477_em-eta17-phi23*/	5,16,3,7,17,3,6,18,1,16,19,1,1,0,2,3,
/* out0478_em-eta18-phi23*/	3,16,0,4,16,3,8,0,2,1,
/* out0479_em-eta19-phi23*/	1,16,0,9
};