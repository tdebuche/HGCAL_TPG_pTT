parameter integer matrixH [0:7637] = {
/* num inputs = 148(in0-in147) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2385 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	3,79,0,2,79,1,3,79,2,1,
/* out0003_em-eta3-phi0*/	5,78,0,15,78,1,8,78,2,11,79,1,4,79,2,3,
/* out0004_em-eta4-phi0*/	4,61,0,8,61,1,2,78,1,2,78,2,5,
/* out0005_em-eta5-phi0*/	3,60,0,9,60,1,13,60,2,2,
/* out0006_em-eta6-phi0*/	3,41,0,2,60,0,7,60,2,3,
/* out0007_em-eta7-phi0*/	2,40,1,6,41,0,1,
/* out0008_em-eta8-phi0*/	2,40,0,12,40,1,4,
/* out0009_em-eta9-phi0*/	4,40,0,4,42,0,16,42,1,5,42,2,1,
/* out0010_em-eta10-phi0*/	3,33,0,3,42,1,2,42,2,12,
/* out0011_em-eta11-phi0*/	6,19,0,14,19,1,10,19,2,3,33,0,10,33,1,3,33,2,2,
/* out0012_em-eta12-phi0*/	8,19,0,2,19,2,6,19,3,16,20,3,6,20,4,2,24,0,2,33,1,1,33,2,13,
/* out0013_em-eta13-phi0*/	4,20,2,1,20,3,7,24,0,11,24,1,1,
/* out0014_em-eta14-phi0*/	3,24,0,1,24,1,1,24,2,10,
/* out0015_em-eta15-phi0*/	2,15,0,4,24,2,3,
/* out0016_em-eta16-phi0*/	3,1,1,6,15,0,6,15,2,1,
/* out0017_em-eta17-phi0*/	3,0,1,11,1,1,2,15,2,5,
/* out0018_em-eta18-phi0*/	3,0,0,7,0,1,4,15,2,3,
/* out0019_em-eta19-phi0*/	1,0,0,6,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	5,62,0,1,62,1,1,79,0,9,79,1,5,79,2,3,
/* out0023_em-eta3-phi1*/	9,61,1,2,62,0,15,62,1,6,62,2,11,78,0,1,78,1,6,79,0,5,79,1,4,79,2,9,
/* out0024_em-eta4-phi1*/	6,42,0,1,43,0,1,61,0,6,61,1,12,61,2,14,62,2,1,
/* out0025_em-eta5-phi1*/	6,42,0,13,42,2,2,60,1,3,60,2,8,61,0,2,61,2,2,
/* out0026_em-eta6-phi1*/	4,41,0,11,41,1,8,42,2,2,60,2,3,
/* out0027_em-eta7-phi1*/	4,22,0,1,40,1,4,41,0,2,41,2,12,
/* out0028_em-eta8-phi1*/	3,22,0,1,40,1,2,40,2,12,
/* out0029_em-eta9-phi1*/	7,21,0,3,21,1,7,40,2,4,42,1,5,43,0,2,50,1,4,50,2,13,
/* out0030_em-eta10-phi1*/	8,19,1,1,20,1,2,21,0,9,33,0,1,42,1,4,42,2,3,43,0,9,43,2,3,
/* out0031_em-eta11-phi1*/	10,19,1,5,19,2,4,19,4,4,19,5,1,20,0,9,20,1,14,33,0,2,33,1,8,34,0,1,43,2,5,
/* out0032_em-eta12-phi1*/	10,19,2,3,20,0,7,20,3,2,20,4,14,20,5,5,24,0,1,33,1,4,33,2,1,34,0,5,34,2,1,
/* out0033_em-eta13-phi1*/	7,2,0,5,20,2,14,20,3,1,20,5,1,24,0,1,24,1,7,34,2,2,
/* out0034_em-eta14-phi1*/	4,2,0,5,2,3,3,24,1,7,24,2,1,
/* out0035_em-eta15-phi1*/	6,0,4,3,2,3,3,15,0,5,15,1,2,24,2,2,25,2,1,
/* out0036_em-eta16-phi1*/	6,0,4,7,1,0,1,1,1,6,15,0,1,15,1,5,15,2,1,
/* out0037_em-eta17-phi1*/	5,0,2,5,1,0,6,1,1,2,15,1,3,15,2,2,
/* out0038_em-eta18-phi1*/	5,0,0,1,0,1,1,0,2,8,0,3,2,15,2,3,
/* out0039_em-eta19-phi1*/	2,0,0,2,0,3,7,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	1,44,2,2,
/* out0043_em-eta3-phi2*/	7,43,0,3,43,1,5,44,0,1,44,1,15,44,2,10,62,1,9,62,2,4,
/* out0044_em-eta4-phi2*/	5,24,1,1,42,1,2,43,0,12,43,1,6,43,2,14,
/* out0045_em-eta5-phi2*/	5,23,1,1,24,0,2,42,0,2,42,1,14,42,2,8,
/* out0046_em-eta6-phi2*/	4,23,0,7,23,1,5,41,1,7,42,2,4,
/* out0047_em-eta7-phi2*/	5,22,0,7,22,1,5,23,0,3,41,1,1,41,2,4,
/* out0048_em-eta8-phi2*/	6,22,0,7,22,1,1,22,2,8,50,1,1,50,2,2,51,0,1,
/* out0049_em-eta9-phi2*/	9,21,1,9,21,2,4,22,2,1,43,0,2,43,1,1,50,1,11,50,2,1,51,0,11,51,2,3,
/* out0050_em-eta10-phi2*/	6,5,1,1,21,0,3,21,2,8,43,0,3,43,1,11,43,2,2,
/* out0051_em-eta11-phi2*/	9,4,1,11,5,1,6,19,4,12,19,5,3,21,0,1,34,0,5,34,1,1,43,1,2,43,2,6,
/* out0052_em-eta12-phi2*/	8,2,1,2,3,1,1,4,0,7,19,5,12,20,5,8,34,0,5,34,1,3,34,2,3,
/* out0053_em-eta13-phi2*/	8,2,0,4,2,1,14,2,2,3,3,1,1,20,2,1,20,5,2,25,0,2,34,2,8,
/* out0054_em-eta14-phi2*/	5,2,0,2,2,2,10,2,3,8,3,4,2,25,0,8,
/* out0055_em-eta15-phi2*/	6,0,4,2,2,3,2,3,3,13,3,4,1,25,0,1,25,2,6,
/* out0056_em-eta16-phi2*/	6,0,4,4,0,5,9,1,0,2,15,1,3,16,1,1,25,2,2,
/* out0057_em-eta17-phi2*/	4,1,0,7,1,4,5,15,1,2,16,1,2,
/* out0058_em-eta18-phi2*/	7,0,2,3,0,3,2,1,3,1,1,4,7,15,1,1,15,2,1,16,1,2,
/* out0059_em-eta19-phi2*/	2,0,3,5,1,3,5,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	3,26,1,5,44,0,1,44,2,3,
/* out0063_em-eta3-phi3*/	9,25,0,2,25,1,14,25,2,1,26,0,4,26,1,7,43,1,1,44,0,14,44,1,1,44,2,1,
/* out0064_em-eta4-phi3*/	6,24,1,12,24,2,1,25,0,14,25,2,1,43,1,4,43,2,2,
/* out0065_em-eta5-phi3*/	4,23,1,3,24,0,14,24,1,3,24,2,8,
/* out0066_em-eta6-phi3*/	4,8,0,1,23,0,3,23,1,7,23,2,12,
/* out0067_em-eta7-phi3*/	5,7,0,4,7,1,3,22,1,6,23,0,3,23,2,3,
/* out0068_em-eta8-phi3*/	6,6,0,3,6,1,1,7,0,2,22,1,4,22,2,6,51,1,1,
/* out0069_em-eta9-phi3*/	7,6,0,11,6,2,1,21,2,2,22,2,1,51,0,4,51,1,10,51,2,7,
/* out0070_em-eta10-phi3*/	9,4,4,16,4,5,4,5,1,2,6,0,1,6,2,2,21,2,2,43,1,2,44,0,10,51,2,5,
/* out0071_em-eta11-phi3*/	8,4,1,4,4,2,11,5,0,14,5,1,7,5,4,2,34,1,2,44,0,4,44,2,8,
/* out0072_em-eta12-phi3*/	9,2,4,1,3,1,3,4,0,9,4,1,1,4,2,5,4,3,12,34,1,8,35,0,2,44,2,1,
/* out0073_em-eta13-phi3*/	11,2,2,1,2,4,5,2,5,1,3,0,8,3,1,11,25,0,2,25,1,2,34,1,2,34,2,2,35,0,2,35,2,1,
/* out0074_em-eta14-phi3*/	6,2,2,2,3,0,8,3,4,11,3,5,1,25,0,3,25,1,5,
/* out0075_em-eta15-phi3*/	6,3,2,11,3,3,3,3,4,2,3,5,2,25,1,2,25,2,5,
/* out0076_em-eta16-phi3*/	6,0,5,7,1,5,6,3,2,2,27,1,1,16,2,3,25,2,2,
/* out0077_em-eta17-phi3*/	5,1,2,1,1,4,2,1,5,9,16,1,3,16,2,1,
/* out0078_em-eta18-phi3*/	4,1,2,5,1,3,4,1,4,2,16,1,3,
/* out0079_em-eta19-phi3*/	3,1,2,1,1,3,6,12,5,4,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	1,26,1,2,
/* out0083_em-eta3-phi4*/	7,10,0,16,10,1,4,10,2,4,25,1,2,25,2,6,26,0,12,26,1,2,
/* out0084_em-eta4-phi4*/	6,9,0,7,9,1,14,9,2,2,10,2,2,24,2,2,25,2,8,
/* out0085_em-eta5-phi4*/	4,8,1,14,8,2,1,9,0,8,24,2,5,
/* out0086_em-eta6-phi4*/	5,7,1,4,8,0,15,8,1,1,8,2,3,23,2,1,
/* out0087_em-eta7-phi4*/	3,7,0,4,7,1,9,7,2,7,
/* out0088_em-eta8-phi4*/	3,6,1,7,7,0,6,7,2,2,
/* out0089_em-eta9-phi4*/	7,6,0,1,6,1,6,6,2,6,51,1,5,52,0,16,52,1,3,52,2,2,
/* out0090_em-eta10-phi4*/	8,4,5,11,5,5,5,6,2,6,63,0,2,44,0,2,44,1,9,51,2,1,52,2,5,
/* out0091_em-eta11-phi4*/	8,4,5,1,5,0,2,5,2,9,5,3,2,5,4,12,5,5,11,44,1,7,44,2,6,
/* out0092_em-eta12-phi4*/	9,4,3,4,5,2,3,5,3,14,5,4,2,45,0,6,45,1,1,35,0,10,35,1,1,44,2,1,
/* out0093_em-eta13-phi4*/	6,2,4,10,2,5,4,45,0,9,45,3,3,35,0,2,35,2,8,
/* out0094_em-eta14-phi4*/	7,2,5,11,3,5,8,27,4,1,45,3,1,25,1,4,26,0,2,35,2,2,
/* out0095_em-eta15-phi4*/	6,3,2,3,3,5,5,27,4,3,28,1,8,25,1,3,26,0,3,
/* out0096_em-eta16-phi4*/	4,27,1,10,28,1,5,16,2,5,26,2,1,
/* out0097_em-eta17-phi4*/	7,1,2,3,1,5,1,27,0,5,27,1,3,16,0,1,16,1,1,16,2,3,
/* out0098_em-eta18-phi4*/	4,1,2,6,12,2,5,27,0,2,16,1,3,
/* out0099_em-eta19-phi4*/	6,11,1,1,11,5,16,12,1,16,12,2,3,12,4,1,12,5,11,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	2,10,1,12,10,2,8,
/* out0104_em-eta4-phi5*/	6,9,1,2,9,2,11,10,2,2,105,1,3,117,1,2,117,2,3,
/* out0105_em-eta5-phi5*/	6,8,1,1,8,2,5,9,0,1,9,2,3,105,0,10,105,1,9,
/* out0106_em-eta6-phi5*/	4,8,2,7,92,0,10,92,1,4,105,0,2,
/* out0107_em-eta7-phi5*/	5,7,2,6,80,0,1,80,1,2,92,0,6,92,2,4,
/* out0108_em-eta8-phi5*/	4,7,2,1,80,0,12,80,1,2,80,2,1,
/* out0109_em-eta9-phi5*/	8,6,1,2,6,2,1,63,0,2,63,1,3,80,0,3,80,2,3,52,1,12,52,2,1,
/* out0110_em-eta10-phi5*/	5,63,0,9,63,1,1,45,0,8,52,1,1,52,2,8,
/* out0111_em-eta11-phi5*/	7,5,2,4,45,1,1,46,1,4,63,0,3,63,2,4,45,0,8,45,2,6,
/* out0112_em-eta12-phi5*/	6,45,1,14,45,2,5,46,0,4,46,1,8,35,1,10,45,2,2,
/* out0113_em-eta13-phi5*/	7,45,0,1,45,2,11,45,3,8,46,3,1,46,4,4,35,1,5,35,2,4,
/* out0114_em-eta14-phi5*/	6,27,4,6,27,5,1,45,3,4,46,3,11,26,0,7,35,2,1,
/* out0115_em-eta15-phi5*/	6,27,4,6,27,5,3,28,0,6,28,1,3,26,0,4,26,2,3,
/* out0116_em-eta16-phi5*/	5,27,1,1,27,2,8,28,0,6,16,2,2,26,2,4,
/* out0117_em-eta17-phi5*/	6,27,0,4,27,1,1,27,2,4,27,3,3,16,0,8,16,2,2,
/* out0118_em-eta18-phi5*/	6,12,2,6,12,3,2,27,0,5,27,3,1,16,0,7,16,1,1,
/* out0119_em-eta19-phi5*/	6,11,1,2,11,2,4,12,2,2,12,3,2,12,4,11,12,5,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	4,117,1,5,129,0,15,129,1,4,129,2,1,
/* out0124_em-eta4-phi6*/	8,105,1,2,105,2,1,117,1,9,117,2,13,118,0,4,118,1,9,129,0,1,129,2,2,
/* out0125_em-eta5-phi6*/	5,105,0,2,105,1,2,105,2,15,106,1,5,118,0,4,
/* out0126_em-eta6-phi6*/	5,92,1,12,92,2,2,105,0,2,106,0,6,106,1,2,
/* out0127_em-eta7-phi6*/	4,80,1,3,92,2,10,93,0,2,93,1,4,
/* out0128_em-eta8-phi6*/	3,80,1,9,80,2,6,93,0,1,
/* out0129_em-eta9-phi6*/	6,63,1,4,80,2,6,81,0,3,53,0,15,53,1,6,53,2,2,
/* out0130_em-eta10-phi6*/	5,63,1,7,63,2,4,45,1,8,53,0,1,53,2,8,
/* out0131_em-eta11-phi6*/	5,45,4,5,63,2,7,64,0,4,45,1,8,45,2,6,
/* out0132_em-eta12-phi6*/	6,45,4,11,45,5,7,46,0,9,46,1,4,36,0,10,45,2,2,
/* out0133_em-eta13-phi6*/	8,45,5,1,46,0,3,46,2,2,46,3,1,46,4,12,46,5,7,36,0,5,36,2,4,
/* out0134_em-eta14-phi6*/	6,27,5,6,28,5,1,46,2,12,46,3,3,26,1,7,36,2,1,
/* out0135_em-eta15-phi6*/	6,27,5,6,28,0,3,28,4,3,28,5,6,26,1,4,26,2,3,
/* out0136_em-eta16-phi6*/	6,27,2,1,28,0,1,28,3,1,28,4,12,17,2,1,26,2,4,
/* out0137_em-eta17-phi6*/	6,27,2,3,27,3,6,28,3,3,28,4,1,17,1,3,17,2,1,
/* out0138_em-eta18-phi6*/	3,12,3,9,27,3,5,17,1,3,
/* out0139_em-eta19-phi6*/	6,11,0,3,11,1,13,11,2,12,11,3,5,12,3,2,12,4,4,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	1,138,2,2,
/* out0143_em-eta3-phi7*/	6,129,1,12,129,2,11,130,0,6,130,1,2,138,1,3,138,2,11,
/* out0144_em-eta4-phi7*/	6,118,0,2,118,1,7,118,2,14,119,0,2,129,2,2,130,0,8,
/* out0145_em-eta5-phi7*/	5,106,1,8,106,2,7,118,0,6,118,2,2,119,0,5,
/* out0146_em-eta6-phi7*/	5,93,1,3,93,2,1,106,0,10,106,1,1,106,2,8,
/* out0147_em-eta7-phi7*/	3,93,0,4,93,1,9,93,2,7,
/* out0148_em-eta8-phi7*/	3,81,0,2,81,1,6,93,0,8,
/* out0149_em-eta9-phi7*/	7,81,0,9,81,1,2,81,2,3,53,1,10,53,2,1,54,0,10,54,1,1,
/* out0150_em-eta10-phi7*/	9,63,1,1,63,2,1,64,1,5,65,1,11,81,0,2,81,2,3,46,0,9,46,1,2,53,2,5,
/* out0151_em-eta11-phi7*/	8,64,0,9,64,1,11,64,2,12,64,3,2,65,0,2,65,1,1,46,0,7,46,2,6,
/* out0152_em-eta12-phi7*/	8,45,5,7,64,0,3,64,2,2,64,3,14,65,3,4,36,0,1,36,1,10,46,2,1,
/* out0153_em-eta13-phi7*/	8,45,5,1,46,2,1,46,5,9,47,0,1,47,1,11,48,1,2,36,1,2,36,2,8,
/* out0154_em-eta14-phi7*/	9,28,5,1,46,2,1,47,0,13,47,1,4,47,2,1,47,3,2,26,1,2,27,0,4,36,2,2,
/* out0155_em-eta15-phi7*/	6,28,2,4,28,5,7,47,0,2,47,3,6,26,1,3,27,0,3,
/* out0156_em-eta16-phi7*/	5,28,2,11,28,3,3,28,5,1,17,2,5,26,2,1,
/* out0157_em-eta17-phi7*/	5,28,3,8,29,0,3,29,1,1,17,1,2,17,2,3,
/* out0158_em-eta18-phi7*/	6,11,3,5,12,3,1,27,3,1,28,3,1,29,0,6,17,1,3,
/* out0159_em-eta19-phi7*/	2,11,0,6,11,3,6,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	4,138,1,2,138,2,3,139,0,1,139,1,3,
/* out0163_em-eta3-phi8*/	8,130,0,1,130,1,14,130,2,2,131,0,1,138,1,11,139,0,15,139,1,3,139,2,2,
/* out0164_em-eta4-phi8*/	5,119,0,1,119,1,12,130,0,1,130,2,14,131,0,6,
/* out0165_em-eta5-phi8*/	4,107,1,3,119,0,8,119,1,3,119,2,14,
/* out0166_em-eta6-phi8*/	4,106,2,1,107,0,7,107,1,13,107,2,2,
/* out0167_em-eta7-phi8*/	3,93,2,7,94,1,6,107,0,6,
/* out0168_em-eta8-phi8*/	6,81,1,4,93,0,1,93,2,1,94,0,6,94,1,4,54,1,1,
/* out0169_em-eta9-phi8*/	7,81,1,4,81,2,7,82,1,2,94,0,1,54,0,6,54,1,9,54,2,8,
/* out0170_em-eta10-phi8*/	9,64,4,16,64,5,2,65,1,4,81,2,3,82,0,1,82,1,1,46,1,10,47,0,2,54,2,5,
/* out0171_em-eta11-phi8*/	8,64,2,2,64,5,7,65,0,14,65,4,11,65,5,4,37,0,2,46,1,4,46,2,8,
/* out0172_em-eta12-phi8*/	9,47,4,3,48,1,1,65,2,9,65,3,12,65,4,5,65,5,1,36,1,2,37,0,8,46,2,1,
/* out0173_em-eta13-phi8*/	11,47,1,1,47,2,1,47,4,3,48,0,7,48,1,13,27,0,2,27,1,2,36,1,2,36,2,1,37,0,2,37,2,2,
/* out0174_em-eta14-phi8*/	6,47,2,13,47,3,1,48,0,3,48,4,5,27,0,5,27,1,3,
/* out0175_em-eta15-phi8*/	6,47,2,1,47,3,7,48,3,9,48,4,2,27,0,2,27,2,5,
/* out0176_em-eta16-phi8*/	6,28,2,1,29,1,6,30,1,7,48,3,1,17,2,4,27,2,2,
/* out0177_em-eta17-phi8*/	6,29,0,1,29,1,9,29,2,2,17,0,7,17,1,1,17,2,2,
/* out0178_em-eta18-phi8*/	4,29,0,5,29,2,2,29,3,4,17,1,3,
/* out0179_em-eta19-phi8*/	3,11,0,7,29,0,1,29,3,6,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	1,139,1,2,
/* out0183_em-eta3-phi9*/	5,131,1,8,139,1,8,139,2,14,140,0,4,140,1,9,
/* out0184_em-eta4-phi9*/	5,119,1,1,120,1,2,131,0,9,131,1,8,131,2,15,
/* out0185_em-eta5-phi9*/	5,107,2,1,119,2,2,120,0,14,120,1,8,120,2,3,
/* out0186_em-eta6-phi9*/	6,107,0,1,107,2,12,108,0,5,108,1,2,120,0,2,120,2,2,
/* out0187_em-eta7-phi9*/	5,94,1,5,94,2,7,107,0,2,107,2,1,108,0,5,
/* out0188_em-eta8-phi9*/	5,94,0,8,94,1,1,94,2,7,54,1,1,55,0,3,
/* out0189_em-eta9-phi9*/	9,82,1,11,82,2,1,94,0,1,47,0,1,47,1,2,54,1,4,54,2,3,55,0,9,55,2,3,
/* out0190_em-eta10-phi9*/	6,64,5,1,82,0,9,82,1,2,47,0,11,47,1,3,47,2,2,
/* out0191_em-eta11-phi9*/	9,64,5,6,65,5,11,66,1,10,67,1,4,82,0,2,37,0,1,37,1,5,47,0,2,47,2,6,
/* out0192_em-eta12-phi9*/	8,47,4,3,65,2,7,66,0,15,66,1,5,66,3,1,37,0,3,37,1,5,37,2,3,
/* out0193_em-eta13-phi9*/	7,47,4,7,47,5,12,48,0,3,66,0,1,66,3,1,27,1,2,37,2,8,
/* out0194_em-eta14-phi9*/	5,48,0,3,48,2,1,48,4,9,48,5,8,27,1,8,
/* out0195_em-eta15-phi9*/	5,29,4,2,48,2,10,48,3,6,27,1,1,27,2,6,
/* out0196_em-eta16-phi9*/	6,29,4,4,30,0,2,30,1,9,17,0,1,18,0,3,27,2,2,
/* out0197_em-eta17-phi9*/	4,29,2,5,30,0,7,17,0,6,18,0,2,
/* out0198_em-eta18-phi9*/	7,29,2,7,29,3,1,30,3,2,30,4,3,17,0,2,17,1,1,18,0,1,
/* out0199_em-eta19-phi9*/	2,29,3,5,30,3,5,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	5,140,1,1,140,2,1,146,0,9,146,1,3,146,2,5,
/* out0203_em-eta3-phi10*/	10,132,1,1,132,2,1,140,0,11,140,1,6,140,2,15,141,0,6,141,2,1,146,0,5,146,1,9,146,2,4,
/* out0204_em-eta4-phi10*/	6,120,1,1,131,2,1,132,0,11,132,1,15,132,2,6,140,0,1,
/* out0205_em-eta5-phi10*/	5,120,1,5,120,2,9,121,0,8,121,1,3,132,0,4,
/* out0206_em-eta6-phi10*/	5,108,0,2,108,1,14,108,2,3,120,2,2,121,0,3,
/* out0207_em-eta7-phi10*/	4,94,2,1,95,1,4,108,0,4,108,2,10,
/* out0208_em-eta8-phi10*/	3,94,2,1,95,0,4,95,1,10,
/* out0209_em-eta9-phi10*/	6,82,2,10,95,0,4,47,1,2,48,0,5,55,0,4,55,2,13,
/* out0210_em-eta10-phi10*/	7,66,4,3,82,0,4,82,2,5,83,1,1,47,1,9,47,2,3,48,0,4,
/* out0211_em-eta11-phi10*/	9,66,1,1,66,2,2,66,4,10,66,5,1,67,0,11,67,1,12,37,1,1,38,0,8,47,2,5,
/* out0212_em-eta12-phi10*/	10,66,2,14,66,3,5,67,0,2,67,3,1,67,4,8,28,1,1,37,1,5,37,2,1,38,0,4,38,2,1,
/* out0213_em-eta13-phi10*/	9,47,5,4,48,5,1,49,1,1,50,1,3,66,3,9,67,3,8,28,0,7,28,1,1,37,2,2,
/* out0214_em-eta14-phi10*/	7,48,2,2,48,5,7,49,0,2,49,1,11,50,1,1,28,0,7,28,2,1,
/* out0215_em-eta15-phi10*/	7,29,4,3,48,2,3,49,0,12,18,0,2,18,1,2,27,2,1,28,2,1,
/* out0216_em-eta16-phi10*/	5,29,4,7,29,5,6,30,0,1,18,0,5,18,1,1,
/* out0217_em-eta17-phi10*/	5,29,5,2,30,0,6,30,4,5,18,0,3,18,2,2,
/* out0218_em-eta18-phi10*/	5,30,2,1,30,3,2,30,4,8,30,5,1,18,2,2,
/* out0219_em-eta19-phi10*/	2,30,2,2,30,3,7,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	3,146,0,2,146,1,1,146,2,3,
/* out0223_em-eta3-phi11*/	5,141,0,10,141,1,16,141,2,11,146,1,3,146,2,4,
/* out0224_em-eta4-phi11*/	5,132,0,1,132,2,9,133,0,5,133,1,16,141,2,4,
/* out0225_em-eta5-phi11*/	4,121,0,2,121,1,13,121,2,9,133,0,3,
/* out0226_em-eta6-phi11*/	5,108,2,2,109,0,4,109,1,8,121,0,3,121,2,7,
/* out0227_em-eta7-phi11*/	4,95,1,1,95,2,4,108,2,1,109,0,12,
/* out0228_em-eta8-phi11*/	3,95,0,4,95,1,1,95,2,12,
/* out0229_em-eta9-phi11*/	5,83,1,9,95,0,4,48,0,5,48,1,12,48,2,1,
/* out0230_em-eta10-phi11*/	5,83,0,6,83,1,6,38,1,3,48,0,2,48,2,11,
/* out0231_em-eta11-phi11*/	9,66,4,3,66,5,15,67,0,3,67,4,1,67,5,7,83,0,2,38,0,3,38,1,9,38,2,2,
/* out0232_em-eta12-phi11*/	7,67,2,11,67,3,3,67,4,7,67,5,9,28,1,1,38,0,1,38,2,9,
/* out0233_em-eta13-phi11*/	6,49,4,8,50,1,9,67,2,5,67,3,4,28,0,1,28,1,9,
/* out0234_em-eta14-phi11*/	6,49,1,3,49,2,8,50,0,8,50,1,3,28,0,1,28,2,7,
/* out0235_em-eta15-phi11*/	6,49,0,2,49,1,1,49,2,8,49,3,8,18,1,4,28,2,3,
/* out0236_em-eta16-phi11*/	3,29,5,6,49,3,8,18,1,5,
/* out0237_em-eta17-phi11*/	3,29,5,2,30,5,11,18,2,5,
/* out0238_em-eta18-phi11*/	3,30,2,7,30,5,4,18,2,3,
/* out0239_em-eta19-phi11*/	1,30,2,6,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	3,147,0,3,147,1,1,147,2,2,
/* out0243_em-eta3-phi12*/	5,142,0,16,142,1,11,142,2,10,147,0,4,147,1,3,
/* out0244_em-eta4-phi12*/	5,133,0,5,133,2,16,134,0,1,134,1,9,142,2,5,
/* out0245_em-eta5-phi12*/	4,122,0,3,122,1,15,122,2,6,133,0,3,
/* out0246_em-eta6-phi12*/	5,109,1,8,109,2,4,110,0,2,122,0,9,122,1,1,
/* out0247_em-eta7-phi12*/	3,96,1,6,109,2,12,110,0,1,
/* out0248_em-eta8-phi12*/	2,96,0,12,96,1,4,
/* out0249_em-eta9-phi12*/	7,83,2,9,96,0,4,39,1,1,48,1,4,48,2,1,49,0,13,49,2,4,
/* out0250_em-eta10-phi12*/	5,83,0,6,83,2,6,39,0,11,39,1,3,48,2,3,
/* out0251_em-eta11-phi12*/	10,68,4,14,68,5,10,69,0,3,69,1,1,83,0,2,29,1,1,38,1,4,38,2,1,39,0,5,39,2,2,
/* out0252_em-eta12-phi12*/	8,68,1,6,68,2,2,68,4,2,69,0,6,69,1,15,29,0,8,29,1,1,38,2,3,
/* out0253_em-eta13-phi12*/	6,49,4,8,49,5,9,68,0,1,68,1,7,28,1,4,29,0,6,
/* out0254_em-eta14-phi12*/	7,49,5,3,50,0,8,50,4,8,50,5,3,19,0,3,19,1,1,28,2,4,
/* out0255_em-eta15-phi12*/	6,50,2,2,50,3,8,50,4,8,50,5,1,18,1,1,19,0,6,
/* out0256_em-eta16-phi12*/	4,31,4,6,50,3,8,18,1,3,19,0,2,
/* out0257_em-eta17-phi12*/	4,31,4,10,32,1,3,9,1,2,18,2,3,
/* out0258_em-eta18-phi12*/	3,32,1,10,9,1,3,18,2,1,
/* out0259_em-eta19-phi12*/	2,31,1,5,32,1,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	4,143,1,2,147,0,5,147,1,3,147,2,9,
/* out0263_em-eta3-phi13*/	10,134,1,1,134,2,1,142,1,5,142,2,1,143,0,15,143,1,12,143,2,4,147,0,4,147,1,9,147,2,5,
/* out0264_em-eta4-phi13*/	6,123,1,1,134,0,11,134,1,6,134,2,15,135,0,1,143,0,1,
/* out0265_em-eta5-phi13*/	5,122,0,1,122,2,10,123,0,2,123,1,13,134,0,4,
/* out0266_em-eta6-phi13*/	5,110,0,3,110,1,14,110,2,2,122,0,3,123,0,2,
/* out0267_em-eta7-phi13*/	3,96,1,4,110,0,10,110,2,4,
/* out0268_em-eta8-phi13*/	3,96,1,2,96,2,12,97,0,2,
/* out0269_em-eta9-phi13*/	6,84,1,10,96,2,4,39,1,1,40,0,6,49,0,3,49,2,12,
/* out0270_em-eta10-phi13*/	8,68,5,1,69,5,2,83,2,1,84,0,4,84,1,5,39,1,11,39,2,4,40,0,1,
/* out0271_em-eta11-phi13*/	9,68,5,5,69,0,4,69,2,4,69,3,1,69,4,9,69,5,14,29,1,3,30,0,1,39,2,9,
/* out0272_em-eta12-phi13*/	8,68,1,2,68,2,14,68,3,5,69,0,3,69,4,7,29,0,1,29,1,8,29,2,2,
/* out0273_em-eta13-phi13*/	8,49,5,3,50,5,1,51,4,5,68,0,14,68,1,1,68,3,1,29,0,1,29,2,9,
/* out0274_em-eta14-phi13*/	7,49,5,1,50,2,2,50,5,11,51,4,5,52,1,3,19,0,1,19,1,7,
/* out0275_em-eta15-phi13*/	7,31,5,2,32,5,1,50,2,12,52,1,3,19,0,3,19,1,1,19,2,2,
/* out0276_em-eta16-phi13*/	6,31,5,13,32,0,1,32,5,1,9,2,1,19,0,1,19,2,4,
/* out0277_em-eta17-phi13*/	5,31,5,1,32,0,11,32,1,1,9,1,4,9,2,3,
/* out0278_em-eta18-phi13*/	5,31,1,2,31,2,4,32,0,3,32,1,1,9,1,3,
/* out0279_em-eta19-phi13*/	2,31,0,5,31,1,8,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	1,144,1,1,
/* out0283_em-eta3-phi14*/	6,135,1,8,143,1,2,143,2,12,144,0,16,144,1,5,144,2,8,
/* out0284_em-eta4-phi14*/	4,123,2,2,135,0,15,135,1,8,135,2,9,
/* out0285_em-eta5-phi14*/	5,111,1,1,123,0,8,123,1,2,123,2,14,124,1,3,
/* out0286_em-eta6-phi14*/	5,110,1,2,110,2,5,111,0,1,111,1,12,123,0,4,
/* out0287_em-eta7-phi14*/	4,97,1,12,110,2,5,111,0,2,111,1,1,
/* out0288_em-eta8-phi14*/	6,97,0,13,97,1,1,97,2,2,40,1,3,41,0,1,41,1,1,
/* out0289_em-eta9-phi14*/	6,84,1,1,84,2,11,97,0,1,40,0,6,40,1,10,40,2,4,
/* out0290_em-eta10-phi14*/	8,70,4,1,84,0,9,84,2,2,30,0,1,30,1,5,39,2,1,40,0,3,40,2,6,
/* out0291_em-eta11-phi14*/	8,69,2,12,69,3,3,70,4,14,71,1,3,84,0,2,30,0,11,30,1,2,30,2,1,
/* out0292_em-eta12-phi14*/	12,51,5,2,52,5,1,68,3,8,69,3,12,70,1,1,71,1,6,20,0,1,20,1,1,29,1,3,29,2,2,30,0,3,30,2,2,
/* out0293_em-eta13-phi14*/	8,51,4,4,51,5,14,52,0,3,52,5,1,68,0,1,68,3,2,20,0,7,29,2,3,
/* out0294_em-eta14-phi14*/	6,51,2,2,51,4,2,52,0,10,52,1,8,19,1,6,20,0,2,
/* out0295_em-eta15-phi14*/	6,32,5,2,51,1,13,51,2,1,52,1,2,19,1,1,19,2,6,
/* out0296_em-eta16-phi14*/	6,32,2,1,32,4,2,32,5,12,9,2,2,10,0,1,19,2,3,
/* out0297_em-eta17-phi14*/	5,31,2,1,32,0,1,32,4,11,9,1,1,9,2,6,
/* out0298_em-eta18-phi14*/	3,31,2,10,31,3,1,9,1,2,
/* out0299_em-eta19-phi14*/	3,31,0,7,31,1,1,31,3,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	3,144,1,3,145,0,2,145,2,3,
/* out0303_em-eta3-phi15*/	7,135,2,1,136,0,2,136,1,14,136,2,1,144,1,7,144,2,8,145,0,11,
/* out0304_em-eta4-phi15*/	5,124,1,5,124,2,8,135,2,6,136,0,14,136,2,1,
/* out0305_em-eta5-phi15*/	4,111,2,3,124,0,14,124,1,8,124,2,4,
/* out0306_em-eta6-phi15*/	4,111,0,7,111,1,2,111,2,13,112,1,1,
/* out0307_em-eta7-phi15*/	4,97,1,3,97,2,4,98,1,7,111,0,6,
/* out0308_em-eta8-phi15*/	8,85,1,3,85,2,1,97,2,10,98,0,1,98,1,1,41,0,3,41,1,1,41,2,3,
/* out0309_em-eta9-phi15*/	10,84,2,2,85,0,1,85,1,11,31,0,4,31,1,4,40,1,3,40,2,4,41,0,11,41,1,13,41,2,11,
/* out0310_em-eta10-phi15*/	9,70,5,10,71,5,12,84,0,1,84,2,1,85,0,2,85,1,1,30,1,5,31,0,10,40,2,2,
/* out0311_em-eta11-phi15*/	8,70,2,4,70,4,1,70,5,6,71,0,15,71,1,4,71,4,7,30,1,4,30,2,9,
/* out0312_em-eta12-phi15*/	10,52,2,1,52,5,3,70,0,4,70,1,15,70,2,5,71,0,1,71,1,3,20,1,7,21,0,1,30,2,4,
/* out0313_em-eta13-phi15*/	8,52,0,1,52,2,5,52,3,1,52,4,8,52,5,11,20,0,4,20,1,3,20,2,3,
/* out0314_em-eta14-phi15*/	7,51,2,11,51,3,1,52,0,2,52,4,8,10,1,1,20,0,2,20,2,4,
/* out0315_em-eta15-phi15*/	7,51,0,11,51,1,3,51,2,2,51,3,2,10,0,4,10,1,2,19,2,1,
/* out0316_em-eta16-phi15*/	4,32,2,12,33,1,1,51,0,2,10,0,6,
/* out0317_em-eta17-phi15*/	5,32,2,2,32,3,9,32,4,2,9,2,4,10,0,2,
/* out0318_em-eta18-phi15*/	5,31,2,1,31,3,7,32,3,2,32,4,1,9,1,1,
/* out0319_em-eta19-phi15*/	3,13,4,7,31,0,4,31,3,4,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	1,145,2,2,
/* out0323_em-eta3-phi16*/	7,136,1,2,136,2,6,137,0,4,137,1,16,137,2,4,145,0,3,145,2,11,
/* out0324_em-eta4-phi16*/	6,124,2,1,125,0,2,125,1,14,125,2,7,136,2,8,137,0,2,
/* out0325_em-eta5-phi16*/	6,112,1,7,112,2,8,124,0,2,124,2,3,125,0,6,125,1,2,
/* out0326_em-eta6-phi16*/	5,98,1,1,98,2,3,112,0,10,112,1,8,112,2,1,
/* out0327_em-eta7-phi16*/	3,98,0,4,98,1,7,98,2,9,
/* out0328_em-eta8-phi16*/	2,85,2,7,98,0,8,
/* out0329_em-eta9-phi16*/	11,85,0,6,85,1,1,85,2,6,31,1,12,31,2,1,32,0,8,32,1,5,32,2,3,41,0,1,41,1,1,41,2,2,
/* out0330_em-eta10-phi16*/	7,71,2,13,71,5,3,72,1,2,85,0,6,21,1,2,31,0,2,31,2,13,
/* out0331_em-eta11-phi16*/	8,70,2,5,70,3,5,71,2,3,71,3,13,71,4,9,71,5,1,21,0,7,21,1,6,
/* out0332_em-eta12-phi16*/	7,54,1,7,70,0,12,70,2,2,70,3,9,20,1,3,21,0,8,21,2,1,
/* out0333_em-eta13-phi16*/	8,52,2,10,52,3,4,53,0,1,53,1,9,54,1,1,11,0,2,20,1,2,20,2,6,
/* out0334_em-eta14-phi16*/	7,33,4,1,51,3,8,52,3,11,53,0,1,10,1,3,11,0,1,20,2,3,
/* out0335_em-eta15-phi16*/	5,33,4,3,34,1,8,51,0,3,51,3,5,10,1,6,
/* out0336_em-eta16-phi16*/	4,33,1,10,34,1,5,10,0,2,10,2,3,
/* out0337_em-eta17-phi16*/	6,32,2,1,32,3,3,33,0,5,33,1,3,10,0,1,10,2,2,
/* out0338_em-eta18-phi16*/	5,13,5,5,14,5,1,31,3,3,32,3,2,33,0,2,
/* out0339_em-eta19-phi16*/	2,13,4,6,13,5,6,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	2,137,0,8,137,2,12,
/* out0344_em-eta4-phi17*/	5,113,1,3,125,0,4,125,2,9,126,2,5,137,0,2,
/* out0345_em-eta5-phi17*/	4,112,2,5,113,0,10,113,1,9,125,0,4,
/* out0346_em-eta6-phi17*/	5,99,0,2,99,1,12,112,0,6,112,2,2,113,0,2,
/* out0347_em-eta7-phi17*/	5,86,1,1,86,2,2,98,0,2,98,2,4,99,0,10,
/* out0348_em-eta8-phi17*/	4,86,0,1,86,1,12,86,2,2,98,0,1,
/* out0349_em-eta9-phi17*/	12,72,1,2,72,2,3,85,0,1,85,2,2,86,0,3,86,1,3,22,0,2,22,1,7,31,2,1,32,0,8,32,1,11,32,2,13,
/* out0350_em-eta10-phi17*/	6,72,1,9,72,2,1,21,1,1,22,0,13,22,1,1,31,2,1,
/* out0351_em-eta11-phi17*/	8,53,4,5,70,3,1,71,3,3,72,0,4,72,1,3,21,1,7,21,2,6,22,0,1,
/* out0352_em-eta12-phi17*/	7,53,4,11,53,5,4,54,0,9,54,1,7,70,3,1,11,1,3,21,2,9,
/* out0353_em-eta13-phi17*/	8,53,0,2,53,1,7,53,2,12,53,3,1,54,0,3,54,1,1,11,0,5,11,1,5,
/* out0354_em-eta14-phi17*/	6,33,4,6,33,5,1,53,0,12,53,3,3,10,1,1,11,0,7,
/* out0355_em-eta15-phi17*/	7,33,4,6,33,5,3,34,0,6,34,1,3,10,1,3,10,2,3,11,0,1,
/* out0356_em-eta16-phi17*/	4,33,1,1,33,2,8,34,0,6,10,2,6,
/* out0357_em-eta17-phi17*/	5,33,0,4,33,1,1,33,2,4,33,3,3,10,2,2,
/* out0358_em-eta18-phi17*/	3,14,5,9,33,0,5,33,3,1,
/* out0359_em-eta19-phi17*/	6,13,4,3,13,5,5,14,0,12,14,1,13,14,4,4,14,5,2,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	5,126,1,4,126,2,2,127,0,1,127,1,15,127,2,4,
/* out0364_em-eta4-phi18*/	8,113,1,2,113,2,1,114,1,11,114,2,2,126,1,12,126,2,9,127,0,2,127,1,1,
/* out0365_em-eta5-phi18*/	7,100,1,5,100,2,1,113,0,2,113,1,2,113,2,15,114,0,1,114,1,3,
/* out0366_em-eta6-phi18*/	4,99,1,4,99,2,10,100,1,7,113,0,2,
/* out0367_em-eta7-phi18*/	4,86,2,3,87,1,6,99,0,4,99,2,6,
/* out0368_em-eta8-phi18*/	3,86,0,6,86,2,9,87,1,1,
/* out0369_em-eta9-phi18*/	9,72,2,4,73,1,3,86,0,6,13,0,1,22,1,7,22,2,2,23,0,13,23,1,11,23,2,8,
/* out0370_em-eta10-phi18*/	6,72,0,4,72,2,7,12,1,1,13,0,1,22,1,1,22,2,13,
/* out0371_em-eta11-phi18*/	7,53,5,4,54,5,1,55,4,4,72,0,7,12,0,6,12,1,7,22,2,1,
/* out0372_em-eta12-phi18*/	6,53,5,8,54,0,4,54,4,5,54,5,14,11,1,3,12,0,9,
/* out0373_em-eta13-phi18*/	7,53,2,4,53,3,1,54,2,1,54,3,8,54,4,11,11,1,5,11,2,5,
/* out0374_em-eta14-phi18*/	6,33,5,6,34,5,1,53,3,11,54,3,4,5,1,1,11,2,7,
/* out0375_em-eta15-phi18*/	7,33,5,6,34,0,3,34,4,3,34,5,6,5,0,3,5,1,3,11,2,1,
/* out0376_em-eta16-phi18*/	5,33,2,1,34,0,1,34,3,1,34,4,12,5,0,6,
/* out0377_em-eta17-phi18*/	5,33,2,3,33,3,6,34,3,3,34,4,1,5,0,2,
/* out0378_em-eta18-phi18*/	3,14,2,6,14,5,2,33,3,5,
/* out0379_em-eta19-phi18*/	6,14,0,4,14,1,2,14,2,2,14,3,1,14,4,11,14,5,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	1,128,0,2,
/* out0383_em-eta3-phi19*/	6,115,1,6,115,2,2,127,0,11,127,2,12,128,0,11,128,2,3,
/* out0384_em-eta4-phi19*/	6,101,1,1,114,0,7,114,1,2,114,2,14,115,1,8,127,0,2,
/* out0385_em-eta5-phi19*/	5,100,1,1,100,2,14,101,0,2,101,1,3,114,0,8,
/* out0386_em-eta6-phi19*/	4,87,2,4,100,0,15,100,1,3,100,2,1,
/* out0387_em-eta7-phi19*/	3,87,0,4,87,1,7,87,2,9,
/* out0388_em-eta8-phi19*/	4,73,1,2,73,2,6,87,0,6,87,1,2,
/* out0389_em-eta9-phi19*/	11,73,0,3,73,1,9,73,2,2,13,0,1,13,1,12,14,0,2,14,1,1,14,2,1,23,0,3,23,1,5,23,2,8,
/* out0390_em-eta10-phi19*/	9,55,5,5,56,5,11,72,0,1,72,2,1,73,0,3,73,1,2,12,1,2,13,0,13,13,2,2,
/* out0391_em-eta11-phi19*/	8,55,4,9,55,5,11,56,0,12,56,1,2,56,4,2,56,5,1,12,1,6,12,2,7,
/* out0392_em-eta12-phi19*/	9,54,2,6,54,5,1,55,1,4,55,4,3,56,0,2,56,1,14,6,1,3,12,0,1,12,2,8,
/* out0393_em-eta13-phi19*/	8,35,4,1,35,5,11,36,5,2,54,2,9,54,3,3,6,0,6,6,1,2,11,2,2,
/* out0394_em-eta14-phi19*/	9,34,5,1,35,4,13,35,5,4,36,0,1,36,1,2,54,3,1,5,1,3,6,0,3,11,2,1,
/* out0395_em-eta15-phi19*/	5,34,2,4,34,5,7,35,4,2,36,1,6,5,1,6,
/* out0396_em-eta16-phi19*/	5,34,2,11,34,3,3,34,5,1,5,0,3,5,2,2,
/* out0397_em-eta17-phi19*/	5,15,4,3,15,5,1,34,3,8,5,0,2,5,2,1,
/* out0398_em-eta18-phi19*/	4,14,2,5,15,4,6,33,3,1,34,3,1,
/* out0399_em-eta19-phi19*/	6,13,1,16,13,3,16,14,1,1,14,2,3,14,3,11,14,4,1,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	4,116,0,1,116,1,3,128,0,3,128,2,2,
/* out0403_em-eta3-phi20*/	8,102,1,1,115,0,2,115,1,1,115,2,14,116,0,15,116,1,3,116,2,2,128,2,11,
/* out0404_em-eta4-phi20*/	5,101,1,8,101,2,5,102,1,6,115,0,14,115,1,1,
/* out0405_em-eta5-phi20*/	4,88,1,3,101,0,14,101,1,4,101,2,8,
/* out0406_em-eta6-phi20*/	4,88,0,7,88,1,13,88,2,2,100,0,1,
/* out0407_em-eta7-phi20*/	5,74,1,4,74,2,3,87,0,4,87,2,3,88,0,6,
/* out0408_em-eta8-phi20*/	6,73,2,4,74,1,10,87,0,2,14,0,3,14,1,1,14,2,3,
/* out0409_em-eta9-phi20*/	10,57,1,2,73,0,7,73,2,4,8,0,4,8,1,3,13,1,4,13,2,4,14,0,11,14,1,13,14,2,11,
/* out0410_em-eta10-phi20*/	9,56,2,16,56,3,3,56,5,4,57,0,1,57,1,1,73,0,3,7,1,5,8,0,2,13,2,10,
/* out0411_em-eta11-phi20*/	7,55,2,11,55,3,4,56,0,2,56,3,6,56,4,14,7,0,9,7,1,4,
/* out0412_em-eta12-phi20*/	9,36,2,3,36,5,1,55,0,9,55,1,12,55,2,5,55,3,1,6,1,7,7,0,4,12,2,1,
/* out0413_em-eta13-phi20*/	8,35,5,1,36,0,1,36,2,3,36,4,7,36,5,13,6,0,3,6,1,3,6,2,4,
/* out0414_em-eta14-phi20*/	7,35,2,5,36,0,13,36,1,1,36,4,3,5,1,1,6,0,4,6,2,2,
/* out0415_em-eta15-phi20*/	7,35,1,9,35,2,2,36,0,1,36,1,7,1,0,1,5,1,2,5,2,4,
/* out0416_em-eta16-phi20*/	5,15,5,6,16,5,7,34,2,1,35,1,1,5,2,6,
/* out0417_em-eta17-phi20*/	5,15,4,1,15,5,9,16,0,2,0,1,4,5,2,2,
/* out0418_em-eta18-phi20*/	4,15,4,5,16,0,2,16,1,4,0,1,1,
/* out0419_em-eta19-phi20*/	3,14,3,4,15,4,1,16,1,6,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	1,116,1,2,
/* out0423_em-eta3-phi21*/	5,102,2,8,103,1,12,103,2,2,116,1,8,116,2,14,
/* out0424_em-eta4-phi21*/	4,89,1,2,102,0,15,102,1,9,102,2,8,
/* out0425_em-eta5-phi21*/	5,88,2,1,89,0,8,89,1,14,89,2,2,101,2,3,
/* out0426_em-eta6-phi21*/	5,75,1,5,75,2,2,88,0,1,88,2,12,89,0,4,
/* out0427_em-eta7-phi21*/	4,74,2,12,75,1,5,88,0,2,88,2,1,
/* out0428_em-eta8-phi21*/	6,74,0,13,74,1,2,74,2,1,8,1,3,14,1,1,14,2,1,
/* out0429_em-eta9-phi21*/	6,57,1,11,57,2,1,74,0,1,8,0,4,8,1,10,8,2,6,
/* out0430_em-eta10-phi21*/	8,56,3,1,57,0,9,57,1,2,3,0,1,7,1,5,7,2,1,8,0,6,8,2,3,
/* out0431_em-eta11-phi21*/	8,37,4,12,38,1,3,55,3,11,56,3,6,57,0,2,7,0,1,7,1,2,7,2,11,
/* out0432_em-eta12-phi21*/	10,36,2,3,37,1,8,38,1,12,55,0,7,2,0,2,2,1,3,6,1,1,6,2,1,7,0,2,7,2,3,
/* out0433_em-eta13-phi21*/	7,36,2,7,36,3,12,36,4,3,37,0,1,37,1,2,2,0,3,6,2,7,
/* out0434_em-eta14-phi21*/	6,35,0,1,35,2,9,35,3,8,36,4,3,1,1,6,6,2,2,
/* out0435_em-eta15-phi21*/	5,16,2,2,35,0,10,35,1,6,1,0,6,1,1,1,
/* out0436_em-eta16-phi21*/	7,16,2,4,16,4,2,16,5,9,0,1,1,0,2,2,1,0,3,5,2,1,
/* out0437_em-eta17-phi21*/	4,16,0,5,16,4,7,0,1,5,0,2,2,
/* out0438_em-eta18-phi21*/	5,15,1,2,15,2,3,16,0,7,16,1,1,0,1,2,
/* out0439_em-eta19-phi21*/	2,15,1,5,16,1,5,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	4,103,2,2,104,0,3,104,1,5,104,2,9,
/* out0443_em-eta3-phi22*/	10,90,1,1,90,2,1,91,0,6,91,2,1,103,0,15,103,1,4,103,2,12,104,0,9,104,1,4,104,2,5,
/* out0444_em-eta4-phi22*/	6,89,2,1,90,0,11,90,1,15,90,2,6,102,0,1,103,0,1,
/* out0445_em-eta5-phi22*/	5,76,0,1,76,1,10,89,0,2,89,2,13,90,0,4,
/* out0446_em-eta6-phi22*/	5,75,0,3,75,1,2,75,2,14,76,0,3,89,0,2,
/* out0447_em-eta7-phi22*/	3,58,2,4,75,0,10,75,1,4,
/* out0448_em-eta8-phi22*/	3,58,1,12,58,2,2,74,0,2,
/* out0449_em-eta9-phi22*/	6,57,2,10,58,1,4,3,1,1,4,0,12,4,2,3,8,2,6,
/* out0450_em-eta10-phi22*/	9,37,5,2,38,5,1,39,0,7,39,1,1,57,0,4,57,2,5,3,0,4,3,1,11,8,2,1,
/* out0451_em-eta11-phi22*/	9,37,4,4,37,5,14,38,0,9,38,1,1,38,4,4,38,5,5,2,1,3,3,0,9,7,2,1,
/* out0452_em-eta12-phi22*/	8,37,1,5,37,2,14,37,3,2,38,0,7,38,4,3,2,0,2,2,1,8,2,2,1,
/* out0453_em-eta13-phi22*/	9,17,5,1,18,5,3,35,3,1,36,3,4,37,0,14,37,1,1,37,3,1,2,0,9,2,2,1,
/* out0454_em-eta14-phi22*/	7,17,4,2,17,5,11,18,5,1,35,0,2,35,3,7,1,1,7,1,2,1,
/* out0455_em-eta15-phi22*/	6,16,2,3,17,4,12,35,0,3,1,0,2,1,1,1,1,2,3,
/* out0456_em-eta16-phi22*/	6,16,2,7,16,3,6,16,4,1,0,2,1,1,0,4,1,2,1,
/* out0457_em-eta17-phi22*/	4,15,2,5,16,3,2,16,4,6,0,2,6,
/* out0458_em-eta18-phi22*/	6,15,0,1,15,1,2,15,2,8,15,3,1,0,1,2,0,2,1,
/* out0459_em-eta19-phi22*/	2,15,0,2,15,1,7,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	3,104,0,1,104,1,3,104,2,2,
/* out0463_em-eta3-phi23*/	5,91,0,10,91,1,16,91,2,11,104,0,3,104,1,4,
/* out0464_em-eta4-phi23*/	5,77,0,5,77,1,16,90,0,1,90,2,9,91,2,4,
/* out0465_em-eta5-phi23*/	4,76,0,3,76,1,6,76,2,15,77,0,11,
/* out0466_em-eta6-phi23*/	5,59,1,4,59,2,8,75,0,2,76,0,9,76,2,1,
/* out0467_em-eta7-phi23*/	4,58,2,6,59,1,12,59,2,8,75,0,1,
/* out0468_em-eta8-phi23*/	2,58,0,12,58,2,4,
/* out0469_em-eta9-phi23*/	6,39,1,9,39,2,1,58,0,4,3,1,1,4,0,4,4,2,13,
/* out0470_em-eta10-phi23*/	5,39,0,6,39,1,6,39,2,15,3,1,3,3,2,11,
/* out0471_em-eta11-phi23*/	8,38,2,14,38,3,1,38,4,3,38,5,10,39,0,3,2,1,1,3,0,2,3,2,5,
/* out0472_em-eta12-phi23*/	7,37,2,2,37,3,6,38,2,2,38,3,15,38,4,6,2,1,1,2,2,8,
/* out0473_em-eta13-phi23*/	6,18,2,16,18,4,8,18,5,9,37,0,1,37,3,7,2,2,6,
/* out0474_em-eta14-phi23*/	6,17,5,3,18,0,8,18,4,8,18,5,3,1,1,1,1,2,3,
/* out0475_em-eta15-phi23*/	5,17,4,2,17,5,1,18,0,8,18,1,8,1,2,6,
/* out0476_em-eta16-phi23*/	4,16,3,6,17,1,16,18,1,8,1,2,2,
/* out0477_em-eta17-phi23*/	3,15,3,11,16,3,2,0,2,2,
/* out0478_em-eta18-phi23*/	4,15,0,7,15,3,4,0,1,1,0,2,2,
/* out0479_em-eta19-phi23*/	1,15,0,6
};