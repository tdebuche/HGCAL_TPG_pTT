parameter integer matrixH [0:2426] = {
/* num inputs = 166(in0-in165) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 6 */
//* total number of input in adders 973 */

/* out0000_had-eta0-phi0*/	1, 121, 2, 
/* out0001_had-eta1-phi0*/	1, 121, 4, 
/* out0002_had-eta2-phi0*/	2, 120, 3, 121, 2, 
/* out0003_had-eta3-phi0*/	3, 116, 1, 117, 12, 120, 4, 
/* out0004_had-eta4-phi0*/	5, 114, 3, 116, 14, 117, 1, 119, 3, 120, 1, 
/* out0005_had-eta5-phi0*/	3, 113, 9, 116, 1, 119, 4, 
/* out0006_had-eta6-phi0*/	5, 72, 1, 112, 9, 113, 2, 118, 3, 119, 1, 
/* out0007_had-eta7-phi0*/	3, 71, 2, 112, 7, 118, 3, 
/* out0008_had-eta8-phi0*/	2, 71, 5, 118, 2, 
/* out0009_had-eta9-phi0*/	2, 70, 7, 71, 1, 
/* out0010_had-eta10-phi0*/	1, 70, 7, 
/* out0011_had-eta11-phi0*/	2, 17, 2, 70, 1, 
/* out0012_had-eta12-phi0*/	1, 17, 2, 
/* out0013_had-eta13-phi0*/	1, 16, 3, 
/* out0014_had-eta14-phi0*/	1, 16, 4, 
/* out0015_had-eta15-phi0*/	1, 16, 3, 
/* out0016_had-eta16-phi0*/	2, 16, 1, 21, 1, 
/* out0017_had-eta17-phi0*/	1, 21, 1, 
/* out0018_had-eta18-phi0*/	1, 21, 1, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	1, 121, 2, 
/* out0021_had-eta1-phi1*/	1, 121, 4, 
/* out0022_had-eta2-phi1*/	3, 115, 1, 120, 3, 121, 2, 
/* out0023_had-eta3-phi1*/	4, 114, 1, 115, 10, 117, 3, 120, 4, 
/* out0024_had-eta4-phi1*/	4, 73, 1, 114, 11, 119, 3, 120, 1, 
/* out0025_had-eta5-phi1*/	4, 73, 5, 113, 4, 114, 1, 119, 4, 
/* out0026_had-eta6-phi1*/	4, 72, 7, 113, 1, 118, 3, 119, 1, 
/* out0027_had-eta7-phi1*/	3, 71, 2, 72, 4, 118, 3, 
/* out0028_had-eta8-phi1*/	3, 71, 5, 83, 1, 118, 2, 
/* out0029_had-eta9-phi1*/	2, 71, 1, 82, 3, 
/* out0030_had-eta10-phi1*/	3, 17, 1, 70, 1, 82, 3, 
/* out0031_had-eta11-phi1*/	1, 17, 3, 
/* out0032_had-eta12-phi1*/	1, 17, 3, 
/* out0033_had-eta13-phi1*/	3, 16, 1, 17, 1, 22, 1, 
/* out0034_had-eta14-phi1*/	2, 16, 2, 22, 1, 
/* out0035_had-eta15-phi1*/	1, 16, 2, 
/* out0036_had-eta16-phi1*/	1, 21, 1, 
/* out0037_had-eta17-phi1*/	1, 21, 1, 
/* out0038_had-eta18-phi1*/	1, 21, 1, 
/* out0039_had-eta19-phi1*/	1, 21, 1, 
/* out0040_had-eta0-phi2*/	1, 125, 2, 
/* out0041_had-eta1-phi2*/	1, 125, 4, 
/* out0042_had-eta2-phi2*/	3, 75, 1, 124, 3, 125, 2, 
/* out0043_had-eta3-phi2*/	4, 74, 4, 75, 7, 115, 5, 124, 4, 
/* out0044_had-eta4-phi2*/	4, 73, 1, 74, 10, 123, 3, 124, 1, 
/* out0045_had-eta5-phi2*/	3, 73, 8, 85, 1, 123, 4, 
/* out0046_had-eta6-phi2*/	5, 72, 3, 73, 1, 84, 4, 122, 3, 123, 1, 
/* out0047_had-eta7-phi2*/	4, 72, 1, 83, 4, 84, 1, 122, 3, 
/* out0048_had-eta8-phi2*/	2, 83, 5, 122, 2, 
/* out0049_had-eta9-phi2*/	1, 82, 4, 
/* out0050_had-eta10-phi2*/	1, 82, 4, 
/* out0051_had-eta11-phi2*/	2, 17, 2, 23, 1, 
/* out0052_had-eta12-phi2*/	2, 17, 2, 23, 1, 
/* out0053_had-eta13-phi2*/	1, 22, 2, 
/* out0054_had-eta14-phi2*/	1, 22, 2, 
/* out0055_had-eta15-phi2*/	2, 21, 1, 22, 1, 
/* out0056_had-eta16-phi2*/	1, 21, 1, 
/* out0057_had-eta17-phi2*/	1, 21, 1, 
/* out0058_had-eta18-phi2*/	1, 21, 1, 
/* out0059_had-eta19-phi2*/	1, 21, 1, 
/* out0060_had-eta0-phi3*/	1, 125, 2, 
/* out0061_had-eta1-phi3*/	1, 125, 4, 
/* out0062_had-eta2-phi3*/	4, 75, 2, 87, 3, 124, 3, 125, 2, 
/* out0063_had-eta3-phi3*/	4, 75, 6, 86, 6, 87, 5, 124, 4, 
/* out0064_had-eta4-phi3*/	5, 74, 2, 85, 5, 86, 5, 123, 3, 124, 1, 
/* out0065_had-eta5-phi3*/	3, 84, 1, 85, 8, 123, 4, 
/* out0066_had-eta6-phi3*/	3, 84, 8, 122, 3, 123, 1, 
/* out0067_had-eta7-phi3*/	4, 83, 3, 84, 2, 94, 2, 122, 3, 
/* out0068_had-eta8-phi3*/	4, 83, 3, 93, 2, 94, 1, 122, 2, 
/* out0069_had-eta9-phi3*/	2, 82, 1, 93, 4, 
/* out0070_had-eta10-phi3*/	3, 23, 2, 82, 1, 93, 1, 
/* out0071_had-eta11-phi3*/	1, 23, 3, 
/* out0072_had-eta12-phi3*/	2, 22, 1, 23, 2, 
/* out0073_had-eta13-phi3*/	1, 22, 2, 
/* out0074_had-eta14-phi3*/	1, 22, 2, 
/* out0075_had-eta15-phi3*/	1, 22, 1, 
/* out0076_had-eta16-phi3*/	1, 21, 1, 
/* out0077_had-eta17-phi3*/	1, 21, 1, 
/* out0078_had-eta18-phi3*/	1, 21, 1, 
/* out0079_had-eta19-phi3*/	2, 0, 1, 21, 1, 
/* out0080_had-eta0-phi4*/	1, 129, 2, 
/* out0081_had-eta1-phi4*/	1, 129, 4, 
/* out0082_had-eta2-phi4*/	3, 87, 2, 128, 3, 129, 2, 
/* out0083_had-eta3-phi4*/	4, 86, 3, 87, 6, 97, 8, 128, 4, 
/* out0084_had-eta4-phi4*/	6, 85, 1, 86, 2, 96, 8, 97, 1, 127, 3, 128, 1, 
/* out0085_had-eta5-phi4*/	4, 85, 1, 95, 6, 96, 2, 127, 4, 
/* out0086_had-eta6-phi4*/	4, 94, 2, 95, 6, 126, 3, 127, 1, 
/* out0087_had-eta7-phi4*/	2, 94, 7, 126, 3, 
/* out0088_had-eta8-phi4*/	3, 93, 3, 94, 2, 126, 2, 
/* out0089_had-eta9-phi4*/	1, 93, 4, 
/* out0090_had-eta10-phi4*/	2, 23, 2, 93, 1, 
/* out0091_had-eta11-phi4*/	1, 23, 3, 
/* out0092_had-eta12-phi4*/	2, 3, 1, 23, 2, 
/* out0093_had-eta13-phi4*/	2, 3, 1, 22, 1, 
/* out0094_had-eta14-phi4*/	1, 22, 2, 
/* out0095_had-eta15-phi4*/	1, 1, 1, 
/* out0096_had-eta16-phi4*/	1, 1, 1, 
/* out0097_had-eta17-phi4*/	1, 1, 1, 
/* out0098_had-eta18-phi4*/	1, 0, 1, 
/* out0099_had-eta19-phi4*/	1, 0, 2, 
/* out0100_had-eta0-phi5*/	1, 129, 2, 
/* out0101_had-eta1-phi5*/	1, 129, 4, 
/* out0102_had-eta2-phi5*/	2, 128, 3, 129, 2, 
/* out0103_had-eta3-phi5*/	2, 97, 7, 128, 4, 
/* out0104_had-eta4-phi5*/	4, 27, 1, 96, 5, 127, 3, 128, 1, 
/* out0105_had-eta5-phi5*/	4, 27, 6, 95, 2, 96, 1, 127, 4, 
/* out0106_had-eta6-phi5*/	4, 26, 5, 95, 2, 126, 3, 127, 1, 
/* out0107_had-eta7-phi5*/	4, 25, 1, 26, 3, 94, 2, 126, 3, 
/* out0108_had-eta8-phi5*/	2, 25, 5, 126, 2, 
/* out0109_had-eta9-phi5*/	3, 24, 2, 25, 2, 93, 1, 
/* out0110_had-eta10-phi5*/	1, 24, 4, 
/* out0111_had-eta11-phi5*/	2, 3, 1, 24, 2, 
/* out0112_had-eta12-phi5*/	1, 3, 2, 
/* out0113_had-eta13-phi5*/	1, 3, 2, 
/* out0114_had-eta14-phi5*/	2, 1, 1, 3, 1, 
/* out0115_had-eta15-phi5*/	1, 1, 2, 
/* out0116_had-eta16-phi5*/	1, 1, 1, 
/* out0117_had-eta17-phi5*/	1, 1, 1, 
/* out0118_had-eta18-phi5*/	1, 0, 2, 
/* out0119_had-eta19-phi5*/	1, 0, 2, 
/* out0120_had-eta0-phi6*/	1, 133, 2, 
/* out0121_had-eta1-phi6*/	1, 133, 4, 
/* out0122_had-eta2-phi6*/	2, 132, 3, 133, 2, 
/* out0123_had-eta3-phi6*/	2, 36, 7, 132, 4, 
/* out0124_had-eta4-phi6*/	4, 27, 2, 35, 5, 131, 3, 132, 1, 
/* out0125_had-eta5-phi6*/	4, 27, 7, 34, 2, 35, 1, 131, 4, 
/* out0126_had-eta6-phi6*/	4, 26, 5, 34, 2, 130, 3, 131, 1, 
/* out0127_had-eta7-phi6*/	4, 25, 1, 26, 3, 33, 2, 130, 3, 
/* out0128_had-eta8-phi6*/	2, 25, 5, 130, 2, 
/* out0129_had-eta9-phi6*/	3, 24, 2, 25, 2, 32, 1, 
/* out0130_had-eta10-phi6*/	1, 24, 4, 
/* out0131_had-eta11-phi6*/	2, 3, 1, 24, 2, 
/* out0132_had-eta12-phi6*/	1, 3, 2, 
/* out0133_had-eta13-phi6*/	1, 3, 2, 
/* out0134_had-eta14-phi6*/	2, 1, 1, 3, 1, 
/* out0135_had-eta15-phi6*/	1, 1, 2, 
/* out0136_had-eta16-phi6*/	1, 1, 1, 
/* out0137_had-eta17-phi6*/	1, 1, 1, 
/* out0138_had-eta18-phi6*/	1, 0, 2, 
/* out0139_had-eta19-phi6*/	1, 0, 2, 
/* out0140_had-eta0-phi7*/	1, 133, 2, 
/* out0141_had-eta1-phi7*/	1, 133, 4, 
/* out0142_had-eta2-phi7*/	3, 47, 2, 132, 3, 133, 2, 
/* out0143_had-eta3-phi7*/	4, 36, 8, 46, 3, 47, 6, 132, 4, 
/* out0144_had-eta4-phi7*/	6, 35, 8, 36, 1, 45, 1, 46, 2, 131, 3, 132, 1, 
/* out0145_had-eta5-phi7*/	4, 34, 6, 35, 2, 45, 1, 131, 4, 
/* out0146_had-eta6-phi7*/	4, 33, 2, 34, 6, 130, 3, 131, 1, 
/* out0147_had-eta7-phi7*/	2, 33, 7, 130, 3, 
/* out0148_had-eta8-phi7*/	3, 32, 3, 33, 2, 130, 2, 
/* out0149_had-eta9-phi7*/	1, 32, 4, 
/* out0150_had-eta10-phi7*/	2, 9, 2, 32, 1, 
/* out0151_had-eta11-phi7*/	1, 9, 3, 
/* out0152_had-eta12-phi7*/	2, 3, 1, 9, 2, 
/* out0153_had-eta13-phi7*/	2, 3, 1, 8, 1, 
/* out0154_had-eta14-phi7*/	1, 8, 2, 
/* out0155_had-eta15-phi7*/	1, 1, 1, 
/* out0156_had-eta16-phi7*/	1, 1, 1, 
/* out0157_had-eta17-phi7*/	1, 1, 1, 
/* out0158_had-eta18-phi7*/	1, 0, 1, 
/* out0159_had-eta19-phi7*/	1, 0, 2, 
/* out0160_had-eta0-phi8*/	1, 137, 2, 
/* out0161_had-eta1-phi8*/	1, 137, 4, 
/* out0162_had-eta2-phi8*/	4, 47, 3, 58, 2, 136, 3, 137, 2, 
/* out0163_had-eta3-phi8*/	4, 46, 6, 47, 5, 58, 6, 136, 4, 
/* out0164_had-eta4-phi8*/	5, 45, 5, 46, 5, 57, 2, 135, 3, 136, 1, 
/* out0165_had-eta5-phi8*/	3, 44, 1, 45, 8, 135, 4, 
/* out0166_had-eta6-phi8*/	3, 44, 8, 134, 3, 135, 1, 
/* out0167_had-eta7-phi8*/	4, 33, 2, 43, 3, 44, 2, 134, 3, 
/* out0168_had-eta8-phi8*/	4, 32, 2, 33, 1, 43, 3, 134, 2, 
/* out0169_had-eta9-phi8*/	2, 32, 4, 42, 1, 
/* out0170_had-eta10-phi8*/	3, 9, 2, 32, 1, 42, 1, 
/* out0171_had-eta11-phi8*/	1, 9, 3, 
/* out0172_had-eta12-phi8*/	2, 8, 1, 9, 2, 
/* out0173_had-eta13-phi8*/	1, 8, 2, 
/* out0174_had-eta14-phi8*/	1, 8, 2, 
/* out0175_had-eta15-phi8*/	1, 8, 1, 
/* out0176_had-eta16-phi8*/	1, 2, 1, 
/* out0177_had-eta17-phi8*/	1, 2, 1, 
/* out0178_had-eta18-phi8*/	1, 2, 1, 
/* out0179_had-eta19-phi8*/	2, 0, 1, 2, 1, 
/* out0180_had-eta0-phi9*/	1, 137, 2, 
/* out0181_had-eta1-phi9*/	1, 137, 4, 
/* out0182_had-eta2-phi9*/	3, 58, 1, 136, 3, 137, 2, 
/* out0183_had-eta3-phi9*/	4, 57, 4, 58, 7, 100, 5, 136, 4, 
/* out0184_had-eta4-phi9*/	4, 56, 1, 57, 10, 135, 3, 136, 1, 
/* out0185_had-eta5-phi9*/	3, 45, 1, 56, 8, 135, 4, 
/* out0186_had-eta6-phi9*/	5, 44, 4, 55, 3, 56, 1, 134, 3, 135, 1, 
/* out0187_had-eta7-phi9*/	4, 43, 4, 44, 1, 55, 1, 134, 3, 
/* out0188_had-eta8-phi9*/	2, 43, 5, 134, 2, 
/* out0189_had-eta9-phi9*/	1, 42, 4, 
/* out0190_had-eta10-phi9*/	1, 42, 4, 
/* out0191_had-eta11-phi9*/	2, 9, 1, 10, 2, 
/* out0192_had-eta12-phi9*/	2, 9, 1, 10, 2, 
/* out0193_had-eta13-phi9*/	1, 8, 2, 
/* out0194_had-eta14-phi9*/	1, 8, 2, 
/* out0195_had-eta15-phi9*/	2, 2, 1, 8, 1, 
/* out0196_had-eta16-phi9*/	1, 2, 1, 
/* out0197_had-eta17-phi9*/	1, 2, 1, 
/* out0198_had-eta18-phi9*/	1, 2, 1, 
/* out0199_had-eta19-phi9*/	1, 2, 1, 
/* out0200_had-eta0-phi10*/	1, 141, 2, 
/* out0201_had-eta1-phi10*/	1, 141, 4, 
/* out0202_had-eta2-phi10*/	3, 100, 1, 140, 3, 141, 2, 
/* out0203_had-eta3-phi10*/	4, 99, 1, 100, 10, 101, 3, 140, 4, 
/* out0204_had-eta4-phi10*/	4, 56, 1, 99, 11, 139, 3, 140, 1, 
/* out0205_had-eta5-phi10*/	4, 56, 5, 98, 4, 99, 1, 139, 4, 
/* out0206_had-eta6-phi10*/	4, 55, 7, 98, 1, 138, 3, 139, 1, 
/* out0207_had-eta7-phi10*/	3, 54, 2, 55, 4, 138, 3, 
/* out0208_had-eta8-phi10*/	3, 43, 1, 54, 5, 138, 2, 
/* out0209_had-eta9-phi10*/	2, 42, 3, 54, 1, 
/* out0210_had-eta10-phi10*/	2, 10, 1, 42, 3, 
/* out0211_had-eta11-phi10*/	1, 10, 3, 
/* out0212_had-eta12-phi10*/	1, 10, 3, 
/* out0213_had-eta13-phi10*/	2, 8, 1, 10, 1, 
/* out0214_had-eta14-phi10*/	2, 8, 1, 14, 1, 
/* out0215_had-eta15-phi10*/	1, 14, 1, 
/* out0216_had-eta16-phi10*/	1, 2, 1, 
/* out0217_had-eta17-phi10*/	1, 2, 1, 
/* out0218_had-eta18-phi10*/	1, 2, 1, 
/* out0219_had-eta19-phi10*/	1, 2, 1, 
/* out0220_had-eta0-phi11*/	1, 141, 2, 
/* out0221_had-eta1-phi11*/	1, 141, 4, 
/* out0222_had-eta2-phi11*/	2, 140, 3, 141, 2, 
/* out0223_had-eta3-phi11*/	2, 101, 12, 140, 4, 
/* out0224_had-eta4-phi11*/	5, 99, 3, 101, 1, 108, 7, 139, 3, 140, 1, 
/* out0225_had-eta5-phi11*/	3, 98, 9, 108, 1, 139, 4, 
/* out0226_had-eta6-phi11*/	5, 55, 1, 98, 2, 106, 4, 138, 3, 139, 1, 
/* out0227_had-eta7-phi11*/	3, 54, 2, 106, 4, 138, 3, 
/* out0228_had-eta8-phi11*/	2, 54, 5, 138, 2, 
/* out0229_had-eta9-phi11*/	2, 54, 1, 64, 3, 
/* out0230_had-eta10-phi11*/	1, 64, 4, 
/* out0231_had-eta11-phi11*/	1, 10, 2, 
/* out0232_had-eta12-phi11*/	1, 10, 2, 
/* out0233_had-eta13-phi11*/	1, 14, 2, 
/* out0234_had-eta14-phi11*/	1, 14, 2, 
/* out0235_had-eta15-phi11*/	1, 14, 1, 
/* out0236_had-eta16-phi11*/	1, 2, 1, 
/* out0237_had-eta17-phi11*/	1, 2, 1, 
/* out0238_had-eta18-phi11*/	1, 2, 1, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	1, 145, 2, 
/* out0241_had-eta1-phi12*/	1, 145, 4, 
/* out0242_had-eta2-phi12*/	2, 144, 3, 145, 2, 
/* out0243_had-eta3-phi12*/	2, 110, 12, 144, 4, 
/* out0244_had-eta4-phi12*/	5, 108, 7, 109, 3, 110, 1, 143, 3, 144, 1, 
/* out0245_had-eta5-phi12*/	3, 107, 9, 108, 1, 143, 4, 
/* out0246_had-eta6-phi12*/	5, 66, 1, 106, 4, 107, 2, 142, 3, 143, 1, 
/* out0247_had-eta7-phi12*/	3, 65, 2, 106, 4, 142, 3, 
/* out0248_had-eta8-phi12*/	2, 65, 5, 142, 2, 
/* out0249_had-eta9-phi12*/	2, 64, 4, 65, 1, 
/* out0250_had-eta10-phi12*/	1, 64, 4, 
/* out0251_had-eta11-phi12*/	2, 15, 2, 64, 1, 
/* out0252_had-eta12-phi12*/	1, 15, 2, 
/* out0253_had-eta13-phi12*/	1, 14, 2, 
/* out0254_had-eta14-phi12*/	1, 14, 2, 
/* out0255_had-eta15-phi12*/	1, 14, 1, 
/* out0256_had-eta16-phi12*/	2, 14, 1, 18, 1, 
/* out0257_had-eta17-phi12*/	1, 18, 1, 
/* out0258_had-eta18-phi12*/	1, 18, 1, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	1, 145, 2, 
/* out0261_had-eta1-phi13*/	1, 145, 4, 
/* out0262_had-eta2-phi13*/	3, 111, 1, 144, 3, 145, 2, 
/* out0263_had-eta3-phi13*/	4, 109, 1, 110, 3, 111, 10, 144, 4, 
/* out0264_had-eta4-phi13*/	4, 67, 1, 109, 11, 143, 3, 144, 1, 
/* out0265_had-eta5-phi13*/	4, 67, 5, 107, 4, 109, 1, 143, 4, 
/* out0266_had-eta6-phi13*/	4, 66, 7, 107, 1, 142, 3, 143, 1, 
/* out0267_had-eta7-phi13*/	3, 65, 2, 66, 4, 142, 3, 
/* out0268_had-eta8-phi13*/	3, 65, 5, 77, 1, 142, 2, 
/* out0269_had-eta9-phi13*/	2, 65, 1, 76, 3, 
/* out0270_had-eta10-phi13*/	2, 15, 1, 76, 3, 
/* out0271_had-eta11-phi13*/	1, 15, 3, 
/* out0272_had-eta12-phi13*/	1, 15, 3, 
/* out0273_had-eta13-phi13*/	3, 14, 1, 15, 1, 19, 1, 
/* out0274_had-eta14-phi13*/	2, 14, 1, 19, 1, 
/* out0275_had-eta15-phi13*/	1, 14, 1, 
/* out0276_had-eta16-phi13*/	1, 18, 1, 
/* out0277_had-eta17-phi13*/	1, 18, 1, 
/* out0278_had-eta18-phi13*/	1, 18, 1, 
/* out0279_had-eta19-phi13*/	1, 18, 1, 
/* out0280_had-eta0-phi14*/	1, 149, 2, 
/* out0281_had-eta1-phi14*/	1, 149, 4, 
/* out0282_had-eta2-phi14*/	3, 69, 1, 148, 3, 149, 2, 
/* out0283_had-eta3-phi14*/	4, 68, 4, 69, 7, 111, 5, 148, 4, 
/* out0284_had-eta4-phi14*/	4, 67, 1, 68, 10, 147, 3, 148, 1, 
/* out0285_had-eta5-phi14*/	3, 67, 8, 79, 1, 147, 4, 
/* out0286_had-eta6-phi14*/	5, 66, 3, 67, 1, 78, 4, 146, 3, 147, 1, 
/* out0287_had-eta7-phi14*/	4, 66, 1, 77, 4, 78, 1, 146, 3, 
/* out0288_had-eta8-phi14*/	2, 77, 5, 146, 2, 
/* out0289_had-eta9-phi14*/	1, 76, 4, 
/* out0290_had-eta10-phi14*/	1, 76, 4, 
/* out0291_had-eta11-phi14*/	2, 15, 2, 20, 1, 
/* out0292_had-eta12-phi14*/	2, 15, 2, 20, 1, 
/* out0293_had-eta13-phi14*/	1, 19, 2, 
/* out0294_had-eta14-phi14*/	1, 19, 2, 
/* out0295_had-eta15-phi14*/	2, 18, 1, 19, 1, 
/* out0296_had-eta16-phi14*/	1, 18, 1, 
/* out0297_had-eta17-phi14*/	1, 18, 1, 
/* out0298_had-eta18-phi14*/	1, 18, 1, 
/* out0299_had-eta19-phi14*/	1, 18, 1, 
/* out0300_had-eta0-phi15*/	1, 149, 2, 
/* out0301_had-eta1-phi15*/	1, 149, 4, 
/* out0302_had-eta2-phi15*/	4, 69, 2, 81, 3, 148, 3, 149, 2, 
/* out0303_had-eta3-phi15*/	4, 69, 6, 80, 6, 81, 5, 148, 4, 
/* out0304_had-eta4-phi15*/	5, 68, 2, 79, 5, 80, 5, 147, 3, 148, 1, 
/* out0305_had-eta5-phi15*/	3, 78, 1, 79, 8, 147, 4, 
/* out0306_had-eta6-phi15*/	3, 78, 8, 146, 3, 147, 1, 
/* out0307_had-eta7-phi15*/	4, 77, 3, 78, 2, 89, 2, 146, 3, 
/* out0308_had-eta8-phi15*/	4, 77, 3, 88, 2, 89, 1, 146, 2, 
/* out0309_had-eta9-phi15*/	2, 76, 1, 88, 4, 
/* out0310_had-eta10-phi15*/	3, 20, 2, 76, 1, 88, 1, 
/* out0311_had-eta11-phi15*/	1, 20, 3, 
/* out0312_had-eta12-phi15*/	2, 19, 1, 20, 2, 
/* out0313_had-eta13-phi15*/	1, 19, 2, 
/* out0314_had-eta14-phi15*/	1, 19, 2, 
/* out0315_had-eta15-phi15*/	1, 19, 1, 
/* out0316_had-eta16-phi15*/	1, 18, 1, 
/* out0317_had-eta17-phi15*/	1, 18, 1, 
/* out0318_had-eta18-phi15*/	1, 18, 1, 
/* out0319_had-eta19-phi15*/	2, 4, 1, 18, 1, 
/* out0320_had-eta0-phi16*/	1, 153, 2, 
/* out0321_had-eta1-phi16*/	1, 153, 4, 
/* out0322_had-eta2-phi16*/	3, 81, 2, 152, 3, 153, 2, 
/* out0323_had-eta3-phi16*/	4, 80, 3, 81, 6, 92, 8, 152, 4, 
/* out0324_had-eta4-phi16*/	6, 79, 1, 80, 2, 91, 8, 92, 1, 151, 3, 152, 1, 
/* out0325_had-eta5-phi16*/	4, 79, 1, 90, 6, 91, 2, 151, 4, 
/* out0326_had-eta6-phi16*/	4, 89, 2, 90, 6, 150, 3, 151, 1, 
/* out0327_had-eta7-phi16*/	2, 89, 7, 150, 3, 
/* out0328_had-eta8-phi16*/	3, 88, 3, 89, 2, 150, 2, 
/* out0329_had-eta9-phi16*/	1, 88, 4, 
/* out0330_had-eta10-phi16*/	2, 20, 2, 88, 1, 
/* out0331_had-eta11-phi16*/	1, 20, 3, 
/* out0332_had-eta12-phi16*/	2, 7, 1, 20, 2, 
/* out0333_had-eta13-phi16*/	2, 7, 1, 19, 1, 
/* out0334_had-eta14-phi16*/	1, 19, 2, 
/* out0335_had-eta15-phi16*/	1, 6, 1, 
/* out0336_had-eta16-phi16*/	1, 6, 1, 
/* out0337_had-eta17-phi16*/	1, 6, 1, 
/* out0338_had-eta18-phi16*/	1, 4, 1, 
/* out0339_had-eta19-phi16*/	1, 4, 2, 
/* out0340_had-eta0-phi17*/	1, 153, 2, 
/* out0341_had-eta1-phi17*/	1, 153, 4, 
/* out0342_had-eta2-phi17*/	2, 152, 3, 153, 2, 
/* out0343_had-eta3-phi17*/	2, 92, 7, 152, 4, 
/* out0344_had-eta4-phi17*/	4, 31, 1, 91, 5, 151, 3, 152, 1, 
/* out0345_had-eta5-phi17*/	4, 31, 6, 90, 2, 91, 1, 151, 4, 
/* out0346_had-eta6-phi17*/	4, 30, 5, 90, 2, 150, 3, 151, 1, 
/* out0347_had-eta7-phi17*/	4, 29, 1, 30, 3, 89, 2, 150, 3, 
/* out0348_had-eta8-phi17*/	2, 29, 5, 150, 2, 
/* out0349_had-eta9-phi17*/	3, 28, 2, 29, 2, 88, 1, 
/* out0350_had-eta10-phi17*/	1, 28, 4, 
/* out0351_had-eta11-phi17*/	2, 7, 1, 28, 2, 
/* out0352_had-eta12-phi17*/	1, 7, 2, 
/* out0353_had-eta13-phi17*/	1, 7, 2, 
/* out0354_had-eta14-phi17*/	2, 6, 1, 7, 1, 
/* out0355_had-eta15-phi17*/	1, 6, 2, 
/* out0356_had-eta16-phi17*/	1, 6, 1, 
/* out0357_had-eta17-phi17*/	1, 6, 1, 
/* out0358_had-eta18-phi17*/	1, 4, 2, 
/* out0359_had-eta19-phi17*/	1, 4, 2, 
/* out0360_had-eta0-phi18*/	1, 157, 2, 
/* out0361_had-eta1-phi18*/	1, 157, 4, 
/* out0362_had-eta2-phi18*/	2, 156, 3, 157, 2, 
/* out0363_had-eta3-phi18*/	2, 41, 7, 156, 4, 
/* out0364_had-eta4-phi18*/	4, 31, 2, 40, 5, 155, 3, 156, 1, 
/* out0365_had-eta5-phi18*/	4, 31, 7, 39, 2, 40, 1, 155, 4, 
/* out0366_had-eta6-phi18*/	4, 30, 5, 39, 2, 154, 3, 155, 1, 
/* out0367_had-eta7-phi18*/	4, 29, 1, 30, 3, 38, 2, 154, 3, 
/* out0368_had-eta8-phi18*/	2, 29, 5, 154, 2, 
/* out0369_had-eta9-phi18*/	3, 28, 2, 29, 2, 37, 1, 
/* out0370_had-eta10-phi18*/	1, 28, 4, 
/* out0371_had-eta11-phi18*/	2, 7, 1, 28, 2, 
/* out0372_had-eta12-phi18*/	1, 7, 2, 
/* out0373_had-eta13-phi18*/	1, 7, 2, 
/* out0374_had-eta14-phi18*/	2, 6, 1, 7, 1, 
/* out0375_had-eta15-phi18*/	1, 6, 2, 
/* out0376_had-eta16-phi18*/	1, 6, 1, 
/* out0377_had-eta17-phi18*/	1, 6, 1, 
/* out0378_had-eta18-phi18*/	1, 4, 2, 
/* out0379_had-eta19-phi18*/	1, 4, 2, 
/* out0380_had-eta0-phi19*/	1, 157, 2, 
/* out0381_had-eta1-phi19*/	1, 157, 4, 
/* out0382_had-eta2-phi19*/	3, 53, 2, 156, 3, 157, 2, 
/* out0383_had-eta3-phi19*/	4, 41, 8, 52, 3, 53, 6, 156, 4, 
/* out0384_had-eta4-phi19*/	6, 40, 8, 41, 1, 51, 1, 52, 2, 155, 3, 156, 1, 
/* out0385_had-eta5-phi19*/	4, 39, 6, 40, 2, 51, 1, 155, 4, 
/* out0386_had-eta6-phi19*/	4, 38, 2, 39, 6, 154, 3, 155, 1, 
/* out0387_had-eta7-phi19*/	2, 38, 7, 154, 3, 
/* out0388_had-eta8-phi19*/	3, 37, 3, 38, 2, 154, 2, 
/* out0389_had-eta9-phi19*/	1, 37, 4, 
/* out0390_had-eta10-phi19*/	2, 13, 2, 37, 1, 
/* out0391_had-eta11-phi19*/	1, 13, 3, 
/* out0392_had-eta12-phi19*/	2, 7, 1, 13, 2, 
/* out0393_had-eta13-phi19*/	2, 7, 1, 11, 1, 
/* out0394_had-eta14-phi19*/	1, 11, 2, 
/* out0395_had-eta15-phi19*/	1, 6, 1, 
/* out0396_had-eta16-phi19*/	1, 6, 1, 
/* out0397_had-eta17-phi19*/	1, 6, 1, 
/* out0398_had-eta18-phi19*/	1, 4, 1, 
/* out0399_had-eta19-phi19*/	1, 4, 2, 
/* out0400_had-eta0-phi20*/	1, 161, 2, 
/* out0401_had-eta1-phi20*/	1, 161, 4, 
/* out0402_had-eta2-phi20*/	4, 53, 3, 63, 2, 160, 3, 161, 2, 
/* out0403_had-eta3-phi20*/	4, 52, 6, 53, 5, 63, 6, 160, 4, 
/* out0404_had-eta4-phi20*/	5, 51, 5, 52, 5, 62, 2, 159, 3, 160, 1, 
/* out0405_had-eta5-phi20*/	3, 50, 1, 51, 8, 159, 4, 
/* out0406_had-eta6-phi20*/	3, 50, 8, 158, 3, 159, 1, 
/* out0407_had-eta7-phi20*/	4, 38, 2, 49, 3, 50, 2, 158, 3, 
/* out0408_had-eta8-phi20*/	4, 37, 2, 38, 1, 49, 3, 158, 2, 
/* out0409_had-eta9-phi20*/	2, 37, 4, 48, 1, 
/* out0410_had-eta10-phi20*/	3, 13, 2, 37, 1, 48, 1, 
/* out0411_had-eta11-phi20*/	1, 13, 3, 
/* out0412_had-eta12-phi20*/	2, 11, 1, 13, 2, 
/* out0413_had-eta13-phi20*/	1, 11, 2, 
/* out0414_had-eta14-phi20*/	1, 11, 2, 
/* out0415_had-eta15-phi20*/	1, 11, 1, 
/* out0416_had-eta16-phi20*/	1, 5, 1, 
/* out0417_had-eta17-phi20*/	1, 5, 1, 
/* out0418_had-eta18-phi20*/	1, 5, 1, 
/* out0419_had-eta19-phi20*/	2, 4, 1, 5, 1, 
/* out0420_had-eta0-phi21*/	1, 161, 2, 
/* out0421_had-eta1-phi21*/	1, 161, 4, 
/* out0422_had-eta2-phi21*/	3, 63, 1, 160, 3, 161, 2, 
/* out0423_had-eta3-phi21*/	4, 62, 4, 63, 7, 105, 5, 160, 4, 
/* out0424_had-eta4-phi21*/	4, 61, 1, 62, 10, 159, 3, 160, 1, 
/* out0425_had-eta5-phi21*/	3, 51, 1, 61, 8, 159, 4, 
/* out0426_had-eta6-phi21*/	5, 50, 4, 60, 3, 61, 1, 158, 3, 159, 1, 
/* out0427_had-eta7-phi21*/	4, 49, 4, 50, 1, 60, 1, 158, 3, 
/* out0428_had-eta8-phi21*/	2, 49, 5, 158, 2, 
/* out0429_had-eta9-phi21*/	1, 48, 4, 
/* out0430_had-eta10-phi21*/	1, 48, 4, 
/* out0431_had-eta11-phi21*/	2, 12, 2, 13, 1, 
/* out0432_had-eta12-phi21*/	2, 12, 2, 13, 1, 
/* out0433_had-eta13-phi21*/	1, 11, 2, 
/* out0434_had-eta14-phi21*/	1, 11, 2, 
/* out0435_had-eta15-phi21*/	2, 5, 1, 11, 1, 
/* out0436_had-eta16-phi21*/	1, 5, 1, 
/* out0437_had-eta17-phi21*/	1, 5, 1, 
/* out0438_had-eta18-phi21*/	1, 5, 1, 
/* out0439_had-eta19-phi21*/	1, 5, 1, 
/* out0440_had-eta0-phi22*/	1, 165, 2, 
/* out0441_had-eta1-phi22*/	1, 165, 4, 
/* out0442_had-eta2-phi22*/	3, 105, 1, 164, 3, 165, 2, 
/* out0443_had-eta3-phi22*/	4, 103, 1, 104, 3, 105, 10, 164, 4, 
/* out0444_had-eta4-phi22*/	4, 61, 1, 103, 11, 163, 3, 164, 1, 
/* out0445_had-eta5-phi22*/	4, 61, 5, 102, 4, 103, 1, 163, 4, 
/* out0446_had-eta6-phi22*/	4, 60, 7, 102, 1, 162, 3, 163, 1, 
/* out0447_had-eta7-phi22*/	3, 59, 2, 60, 4, 162, 3, 
/* out0448_had-eta8-phi22*/	3, 49, 1, 59, 5, 162, 2, 
/* out0449_had-eta9-phi22*/	2, 48, 3, 59, 1, 
/* out0450_had-eta10-phi22*/	2, 12, 1, 48, 3, 
/* out0451_had-eta11-phi22*/	1, 12, 3, 
/* out0452_had-eta12-phi22*/	1, 12, 3, 
/* out0453_had-eta13-phi22*/	2, 11, 1, 12, 1, 
/* out0454_had-eta14-phi22*/	1, 11, 1, 
/* out0455_had-eta15-phi22*/	0, 
/* out0456_had-eta16-phi22*/	1, 5, 1, 
/* out0457_had-eta17-phi22*/	1, 5, 1, 
/* out0458_had-eta18-phi22*/	1, 5, 1, 
/* out0459_had-eta19-phi22*/	1, 5, 1, 
/* out0460_had-eta0-phi23*/	1, 165, 2, 
/* out0461_had-eta1-phi23*/	1, 165, 4, 
/* out0462_had-eta2-phi23*/	2, 164, 3, 165, 2, 
/* out0463_had-eta3-phi23*/	2, 104, 12, 164, 4, 
/* out0464_had-eta4-phi23*/	4, 103, 3, 104, 1, 163, 3, 164, 1, 
/* out0465_had-eta5-phi23*/	2, 102, 9, 163, 4, 
/* out0466_had-eta6-phi23*/	4, 60, 1, 102, 2, 162, 3, 163, 1, 
/* out0467_had-eta7-phi23*/	2, 59, 2, 162, 3, 
/* out0468_had-eta8-phi23*/	2, 59, 5, 162, 2, 
/* out0469_had-eta9-phi23*/	1, 59, 1, 
/* out0470_had-eta10-phi23*/	0, 
/* out0471_had-eta11-phi23*/	1, 12, 2, 
/* out0472_had-eta12-phi23*/	1, 12, 2, 
/* out0473_had-eta13-phi23*/	0, 
/* out0474_had-eta14-phi23*/	0, 
/* out0475_had-eta15-phi23*/	0, 
/* out0476_had-eta16-phi23*/	1, 5, 1, 
/* out0477_had-eta17-phi23*/	1, 5, 1, 
/* out0478_had-eta18-phi23*/	1, 5, 1, 
/* out0479_had-eta19-phi23*/	0, 
};