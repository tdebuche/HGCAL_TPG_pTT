parameter integer matrixH [0:4206] = {
/* num inputs = 298(in0-in297) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 8 */
//* total number of input in adders 1823 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	1, 0, 1, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	0, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	0, 
/* out0033_had-eta13-phi1*/	1, 3, 1, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	1, 1, 1, 
/* out0036_had-eta16-phi1*/	1, 1, 1, 
/* out0037_had-eta17-phi1*/	1, 1, 1, 
/* out0038_had-eta18-phi1*/	1, 0, 1, 
/* out0039_had-eta19-phi1*/	1, 0, 2, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	1, 28, 7, 
/* out0045_had-eta5-phi2*/	2, 27, 5, 28, 1, 
/* out0046_had-eta6-phi2*/	2, 26, 2, 27, 3, 
/* out0047_had-eta7-phi2*/	1, 26, 5, 
/* out0048_had-eta8-phi2*/	1, 25, 4, 
/* out0049_had-eta9-phi2*/	2, 25, 4, 193, 2, 
/* out0050_had-eta10-phi2*/	2, 24, 4, 192, 1, 
/* out0051_had-eta11-phi2*/	2, 24, 3, 192, 2, 
/* out0052_had-eta12-phi2*/	2, 3, 2, 24, 1, 
/* out0053_had-eta13-phi2*/	2, 3, 2, 191, 2, 
/* out0054_had-eta14-phi2*/	2, 3, 2, 191, 1, 
/* out0055_had-eta15-phi2*/	2, 1, 2, 190, 1, 
/* out0056_had-eta16-phi2*/	2, 1, 1, 190, 1, 
/* out0057_had-eta17-phi2*/	2, 1, 1, 190, 1, 
/* out0058_had-eta18-phi2*/	2, 0, 1, 1, 1, 
/* out0059_had-eta19-phi2*/	1, 0, 3, 
/* out0060_had-eta0-phi3*/	1, 253, 1, 
/* out0061_had-eta1-phi3*/	1, 253, 5, 
/* out0062_had-eta2-phi3*/	3, 39, 5, 252, 2, 253, 2, 
/* out0063_had-eta3-phi3*/	3, 38, 4, 39, 4, 252, 4, 
/* out0064_had-eta4-phi3*/	5, 28, 7, 37, 2, 38, 4, 251, 3, 252, 2, 
/* out0065_had-eta5-phi3*/	4, 27, 5, 28, 1, 37, 4, 251, 4, 
/* out0066_had-eta6-phi3*/	5, 26, 2, 27, 3, 36, 3, 250, 2, 251, 1, 
/* out0067_had-eta7-phi3*/	4, 26, 6, 35, 1, 36, 1, 250, 3, 
/* out0068_had-eta8-phi3*/	6, 25, 4, 26, 1, 35, 1, 193, 3, 245, 2, 250, 2, 
/* out0069_had-eta9-phi3*/	6, 25, 4, 34, 1, 193, 6, 244, 1, 245, 6, 250, 1, 
/* out0070_had-eta10-phi3*/	4, 24, 4, 192, 3, 193, 2, 244, 5, 
/* out0071_had-eta11-phi3*/	4, 24, 3, 192, 4, 243, 1, 244, 1, 
/* out0072_had-eta12-phi3*/	5, 3, 2, 24, 1, 191, 2, 192, 1, 243, 3, 
/* out0073_had-eta13-phi3*/	3, 3, 3, 191, 3, 243, 1, 
/* out0074_had-eta14-phi3*/	3, 3, 2, 191, 2, 242, 2, 
/* out0075_had-eta15-phi3*/	3, 1, 2, 190, 2, 242, 2, 
/* out0076_had-eta16-phi3*/	2, 1, 1, 190, 2, 
/* out0077_had-eta17-phi3*/	3, 1, 1, 190, 2, 241, 2, 
/* out0078_had-eta18-phi3*/	3, 0, 1, 1, 1, 241, 1, 
/* out0079_had-eta19-phi3*/	1, 0, 3, 
/* out0080_had-eta0-phi4*/	1, 253, 1, 
/* out0081_had-eta1-phi4*/	1, 253, 5, 
/* out0082_had-eta2-phi4*/	5, 39, 4, 51, 1, 52, 11, 252, 2, 253, 2, 
/* out0083_had-eta3-phi4*/	4, 38, 4, 39, 3, 51, 7, 252, 4, 
/* out0084_had-eta4-phi4*/	5, 37, 3, 38, 4, 50, 5, 251, 3, 252, 2, 
/* out0085_had-eta5-phi4*/	4, 36, 1, 37, 7, 49, 2, 251, 4, 
/* out0086_had-eta6-phi4*/	3, 36, 8, 250, 2, 251, 1, 
/* out0087_had-eta7-phi4*/	3, 35, 5, 36, 2, 250, 3, 
/* out0088_had-eta8-phi4*/	5, 35, 6, 189, 6, 239, 1, 245, 3, 250, 2, 
/* out0089_had-eta9-phi4*/	8, 34, 5, 188, 3, 189, 3, 193, 3, 239, 2, 244, 2, 245, 5, 250, 1, 
/* out0090_had-eta10-phi4*/	4, 34, 4, 188, 4, 192, 1, 244, 5, 
/* out0091_had-eta11-phi4*/	5, 9, 3, 187, 1, 192, 3, 243, 2, 244, 2, 
/* out0092_had-eta12-phi4*/	5, 9, 3, 187, 2, 191, 1, 192, 1, 243, 4, 
/* out0093_had-eta13-phi4*/	6, 3, 1, 8, 1, 9, 1, 191, 3, 242, 1, 243, 2, 
/* out0094_had-eta14-phi4*/	5, 3, 1, 8, 1, 186, 1, 191, 2, 242, 3, 
/* out0095_had-eta15-phi4*/	4, 1, 1, 8, 1, 190, 2, 242, 2, 
/* out0096_had-eta16-phi4*/	4, 1, 1, 190, 2, 241, 2, 242, 1, 
/* out0097_had-eta17-phi4*/	3, 1, 1, 190, 1, 241, 3, 
/* out0098_had-eta18-phi4*/	3, 0, 1, 2, 1, 241, 1, 
/* out0099_had-eta19-phi4*/	1, 0, 2, 
/* out0100_had-eta0-phi5*/	1, 257, 1, 
/* out0101_had-eta1-phi5*/	1, 257, 5, 
/* out0102_had-eta2-phi5*/	5, 51, 1, 52, 5, 91, 10, 256, 2, 257, 2, 
/* out0103_had-eta3-phi5*/	5, 50, 1, 51, 7, 90, 6, 91, 2, 256, 4, 
/* out0104_had-eta4-phi5*/	5, 50, 10, 89, 2, 90, 1, 255, 3, 256, 2, 
/* out0105_had-eta5-phi5*/	3, 49, 10, 89, 1, 255, 4, 
/* out0106_had-eta6-phi5*/	5, 36, 1, 48, 5, 49, 3, 254, 2, 255, 1, 
/* out0107_had-eta7-phi5*/	4, 35, 1, 47, 1, 48, 5, 254, 3, 
/* out0108_had-eta8-phi5*/	6, 35, 2, 47, 4, 183, 2, 189, 5, 239, 3, 254, 2, 
/* out0109_had-eta9-phi5*/	7, 34, 3, 47, 1, 183, 2, 188, 4, 189, 2, 239, 6, 254, 1, 
/* out0110_had-eta10-phi5*/	5, 34, 3, 46, 1, 188, 5, 237, 4, 239, 2, 
/* out0111_had-eta11-phi5*/	3, 9, 3, 187, 4, 237, 4, 
/* out0112_had-eta12-phi5*/	5, 9, 3, 187, 4, 236, 1, 237, 1, 243, 2, 
/* out0113_had-eta13-phi5*/	6, 8, 2, 9, 1, 186, 2, 187, 1, 236, 2, 243, 1, 
/* out0114_had-eta14-phi5*/	3, 8, 2, 186, 2, 242, 2, 
/* out0115_had-eta15-phi5*/	4, 8, 2, 186, 1, 190, 1, 242, 2, 
/* out0116_had-eta16-phi5*/	6, 2, 1, 8, 1, 185, 1, 190, 1, 241, 2, 242, 1, 
/* out0117_had-eta17-phi5*/	3, 2, 1, 185, 1, 241, 3, 
/* out0118_had-eta18-phi5*/	1, 2, 1, 
/* out0119_had-eta19-phi5*/	2, 0, 1, 2, 1, 
/* out0120_had-eta0-phi6*/	1, 257, 1, 
/* out0121_had-eta1-phi6*/	1, 257, 5, 
/* out0122_had-eta2-phi6*/	5, 91, 4, 102, 7, 104, 1, 256, 2, 257, 2, 
/* out0123_had-eta3-phi6*/	4, 90, 7, 100, 3, 102, 4, 256, 4, 
/* out0124_had-eta4-phi6*/	5, 89, 9, 90, 2, 100, 2, 255, 3, 256, 2, 
/* out0125_had-eta5-phi6*/	4, 49, 1, 88, 5, 89, 4, 255, 4, 
/* out0126_had-eta6-phi6*/	5, 48, 3, 87, 1, 88, 5, 254, 2, 255, 1, 
/* out0127_had-eta7-phi6*/	4, 47, 1, 48, 3, 87, 3, 254, 3, 
/* out0128_had-eta8-phi6*/	3, 47, 6, 183, 4, 254, 2, 
/* out0129_had-eta9-phi6*/	7, 46, 2, 47, 2, 182, 1, 183, 6, 239, 2, 240, 4, 254, 1, 
/* out0130_had-eta10-phi6*/	4, 46, 4, 182, 5, 237, 3, 240, 2, 
/* out0131_had-eta11-phi6*/	5, 9, 1, 46, 2, 182, 2, 187, 2, 237, 4, 
/* out0132_had-eta12-phi6*/	5, 9, 1, 10, 2, 181, 1, 187, 2, 236, 4, 
/* out0133_had-eta13-phi6*/	4, 8, 1, 10, 1, 186, 3, 236, 3, 
/* out0134_had-eta14-phi6*/	4, 8, 2, 186, 2, 235, 1, 236, 1, 
/* out0135_had-eta15-phi6*/	3, 8, 2, 186, 2, 235, 2, 
/* out0136_had-eta16-phi6*/	3, 2, 1, 185, 2, 235, 1, 
/* out0137_had-eta17-phi6*/	3, 2, 1, 185, 2, 241, 2, 
/* out0138_had-eta18-phi6*/	1, 2, 1, 
/* out0139_had-eta19-phi6*/	1, 2, 1, 
/* out0140_had-eta0-phi7*/	1, 261, 1, 
/* out0141_had-eta1-phi7*/	1, 261, 5, 
/* out0142_had-eta2-phi7*/	5, 102, 3, 103, 4, 104, 15, 260, 2, 261, 2, 
/* out0143_had-eta3-phi7*/	5, 100, 7, 101, 1, 102, 2, 103, 6, 260, 4, 
/* out0144_had-eta4-phi7*/	5, 99, 7, 100, 4, 101, 1, 259, 3, 260, 2, 
/* out0145_had-eta5-phi7*/	4, 88, 3, 98, 2, 99, 6, 259, 4, 
/* out0146_had-eta6-phi7*/	5, 87, 3, 88, 3, 98, 3, 258, 2, 259, 1, 
/* out0147_had-eta7-phi7*/	2, 87, 7, 258, 3, 
/* out0148_had-eta8-phi7*/	6, 47, 1, 86, 4, 87, 1, 183, 1, 184, 2, 258, 2, 
/* out0149_had-eta9-phi7*/	7, 46, 2, 86, 3, 182, 1, 183, 1, 184, 5, 240, 6, 258, 1, 
/* out0150_had-eta10-phi7*/	4, 46, 4, 182, 5, 238, 2, 240, 4, 
/* out0151_had-eta11-phi7*/	5, 10, 2, 46, 1, 181, 2, 182, 2, 238, 4, 
/* out0152_had-eta12-phi7*/	4, 10, 3, 181, 4, 236, 2, 238, 2, 
/* out0153_had-eta13-phi7*/	5, 10, 2, 181, 2, 186, 1, 236, 2, 246, 1, 
/* out0154_had-eta14-phi7*/	6, 8, 1, 14, 1, 175, 1, 186, 1, 235, 2, 236, 1, 
/* out0155_had-eta15-phi7*/	5, 14, 1, 175, 1, 185, 1, 186, 1, 235, 2, 
/* out0156_had-eta16-phi7*/	3, 2, 1, 185, 2, 235, 2, 
/* out0157_had-eta17-phi7*/	3, 2, 1, 185, 2, 235, 1, 
/* out0158_had-eta18-phi7*/	2, 2, 1, 185, 1, 
/* out0159_had-eta19-phi7*/	1, 2, 1, 
/* out0160_had-eta0-phi8*/	1, 261, 1, 
/* out0161_had-eta1-phi8*/	1, 261, 5, 
/* out0162_had-eta2-phi8*/	4, 103, 3, 114, 2, 260, 2, 261, 2, 
/* out0163_had-eta3-phi8*/	4, 101, 7, 103, 3, 114, 6, 260, 4, 
/* out0164_had-eta4-phi8*/	5, 99, 2, 101, 7, 112, 4, 259, 3, 260, 2, 
/* out0165_had-eta5-phi8*/	4, 98, 4, 99, 1, 112, 4, 259, 4, 
/* out0166_had-eta6-phi8*/	4, 98, 7, 122, 1, 258, 2, 259, 1, 
/* out0167_had-eta7-phi8*/	3, 87, 1, 122, 6, 258, 3, 
/* out0168_had-eta8-phi8*/	4, 86, 5, 122, 1, 184, 2, 258, 2, 
/* out0169_had-eta9-phi8*/	5, 86, 4, 139, 1, 184, 7, 248, 4, 258, 1, 
/* out0170_had-eta10-phi8*/	4, 139, 4, 177, 5, 238, 2, 248, 3, 
/* out0171_had-eta11-phi8*/	5, 10, 1, 139, 2, 177, 3, 181, 1, 238, 4, 
/* out0172_had-eta12-phi8*/	4, 10, 3, 181, 4, 238, 2, 246, 2, 
/* out0173_had-eta13-phi8*/	5, 10, 2, 14, 1, 175, 1, 181, 2, 246, 3, 
/* out0174_had-eta14-phi8*/	4, 14, 2, 175, 3, 235, 1, 246, 2, 
/* out0175_had-eta15-phi8*/	3, 14, 2, 175, 2, 235, 2, 
/* out0176_had-eta16-phi8*/	3, 14, 1, 185, 1, 235, 2, 
/* out0177_had-eta17-phi8*/	2, 2, 1, 185, 2, 
/* out0178_had-eta18-phi8*/	2, 2, 1, 185, 1, 
/* out0179_had-eta19-phi8*/	1, 2, 1, 
/* out0180_had-eta0-phi9*/	1, 265, 1, 
/* out0181_had-eta1-phi9*/	1, 265, 5, 
/* out0182_had-eta2-phi9*/	4, 114, 2, 115, 3, 264, 2, 265, 2, 
/* out0183_had-eta3-phi9*/	4, 113, 7, 114, 6, 115, 3, 264, 4, 
/* out0184_had-eta4-phi9*/	5, 112, 4, 113, 7, 124, 2, 263, 3, 264, 2, 
/* out0185_had-eta5-phi9*/	4, 112, 4, 123, 4, 124, 1, 263, 4, 
/* out0186_had-eta6-phi9*/	4, 122, 1, 123, 7, 262, 2, 263, 1, 
/* out0187_had-eta7-phi9*/	3, 122, 6, 141, 1, 262, 3, 
/* out0188_had-eta8-phi9*/	4, 122, 1, 140, 5, 179, 2, 262, 2, 
/* out0189_had-eta9-phi9*/	5, 139, 1, 140, 4, 179, 7, 248, 5, 262, 1, 
/* out0190_had-eta10-phi9*/	4, 139, 4, 177, 5, 247, 2, 248, 4, 
/* out0191_had-eta11-phi9*/	5, 15, 1, 139, 3, 176, 1, 177, 3, 247, 4, 
/* out0192_had-eta12-phi9*/	4, 15, 3, 176, 4, 246, 2, 247, 2, 
/* out0193_had-eta13-phi9*/	5, 14, 1, 15, 2, 175, 1, 176, 2, 246, 3, 
/* out0194_had-eta14-phi9*/	4, 14, 2, 175, 3, 231, 1, 246, 2, 
/* out0195_had-eta15-phi9*/	3, 14, 2, 175, 2, 231, 2, 
/* out0196_had-eta16-phi9*/	3, 14, 1, 170, 1, 231, 2, 
/* out0197_had-eta17-phi9*/	2, 18, 1, 170, 2, 
/* out0198_had-eta18-phi9*/	2, 18, 1, 170, 1, 
/* out0199_had-eta19-phi9*/	1, 18, 1, 
/* out0200_had-eta0-phi10*/	1, 265, 1, 
/* out0201_had-eta1-phi10*/	1, 265, 5, 
/* out0202_had-eta2-phi10*/	5, 115, 4, 116, 15, 126, 3, 264, 2, 265, 2, 
/* out0203_had-eta3-phi10*/	5, 113, 1, 115, 6, 125, 7, 126, 2, 264, 4, 
/* out0204_had-eta4-phi10*/	5, 113, 1, 124, 7, 125, 4, 263, 3, 264, 2, 
/* out0205_had-eta5-phi10*/	4, 123, 2, 124, 6, 142, 3, 263, 4, 
/* out0206_had-eta6-phi10*/	5, 123, 3, 141, 3, 142, 3, 262, 2, 263, 1, 
/* out0207_had-eta7-phi10*/	2, 141, 7, 262, 3, 
/* out0208_had-eta8-phi10*/	6, 61, 1, 140, 4, 141, 1, 179, 2, 180, 1, 262, 2, 
/* out0209_had-eta9-phi10*/	7, 60, 2, 140, 3, 178, 1, 179, 5, 180, 1, 249, 6, 262, 1, 
/* out0210_had-eta10-phi10*/	5, 60, 4, 139, 1, 178, 5, 247, 2, 249, 4, 
/* out0211_had-eta11-phi10*/	5, 15, 2, 60, 1, 176, 2, 178, 2, 247, 4, 
/* out0212_had-eta12-phi10*/	4, 15, 3, 176, 4, 232, 2, 247, 2, 
/* out0213_had-eta13-phi10*/	5, 15, 2, 171, 1, 176, 2, 232, 2, 246, 1, 
/* out0214_had-eta14-phi10*/	6, 14, 1, 19, 1, 171, 1, 175, 1, 231, 2, 232, 1, 
/* out0215_had-eta15-phi10*/	5, 14, 1, 170, 1, 171, 1, 175, 1, 231, 2, 
/* out0216_had-eta16-phi10*/	3, 18, 1, 170, 2, 231, 2, 
/* out0217_had-eta17-phi10*/	3, 18, 1, 170, 2, 231, 1, 
/* out0218_had-eta18-phi10*/	2, 18, 1, 170, 1, 
/* out0219_had-eta19-phi10*/	1, 18, 1, 
/* out0220_had-eta0-phi11*/	1, 269, 1, 
/* out0221_had-eta1-phi11*/	1, 269, 5, 
/* out0222_had-eta2-phi11*/	5, 116, 1, 126, 7, 145, 4, 268, 2, 269, 2, 
/* out0223_had-eta3-phi11*/	4, 125, 3, 126, 4, 144, 7, 268, 4, 
/* out0224_had-eta4-phi11*/	5, 125, 2, 143, 9, 144, 2, 267, 3, 268, 2, 
/* out0225_had-eta5-phi11*/	4, 63, 1, 142, 5, 143, 4, 267, 4, 
/* out0226_had-eta6-phi11*/	5, 62, 3, 141, 1, 142, 5, 266, 2, 267, 1, 
/* out0227_had-eta7-phi11*/	4, 61, 1, 62, 3, 141, 3, 266, 3, 
/* out0228_had-eta8-phi11*/	3, 61, 6, 180, 4, 266, 2, 
/* out0229_had-eta9-phi11*/	7, 60, 2, 61, 2, 178, 1, 180, 6, 234, 2, 249, 4, 266, 1, 
/* out0230_had-eta10-phi11*/	4, 60, 4, 178, 5, 233, 3, 249, 2, 
/* out0231_had-eta11-phi11*/	5, 20, 1, 60, 2, 172, 2, 178, 2, 233, 4, 
/* out0232_had-eta12-phi11*/	5, 15, 2, 20, 1, 172, 2, 176, 1, 232, 4, 
/* out0233_had-eta13-phi11*/	4, 15, 1, 19, 1, 171, 3, 232, 3, 
/* out0234_had-eta14-phi11*/	4, 19, 2, 171, 2, 231, 1, 232, 1, 
/* out0235_had-eta15-phi11*/	3, 19, 2, 171, 2, 231, 2, 
/* out0236_had-eta16-phi11*/	3, 18, 1, 170, 2, 231, 1, 
/* out0237_had-eta17-phi11*/	3, 18, 1, 170, 2, 226, 2, 
/* out0238_had-eta18-phi11*/	1, 18, 1, 
/* out0239_had-eta19-phi11*/	1, 18, 1, 
/* out0240_had-eta0-phi12*/	1, 269, 1, 
/* out0241_had-eta1-phi12*/	1, 269, 5, 
/* out0242_had-eta2-phi12*/	5, 65, 1, 66, 5, 145, 10, 268, 2, 269, 2, 
/* out0243_had-eta3-phi12*/	5, 64, 1, 65, 7, 144, 6, 145, 2, 268, 4, 
/* out0244_had-eta4-phi12*/	5, 64, 10, 143, 2, 144, 1, 267, 3, 268, 2, 
/* out0245_had-eta5-phi12*/	3, 63, 10, 143, 1, 267, 4, 
/* out0246_had-eta6-phi12*/	5, 62, 5, 63, 3, 76, 1, 266, 2, 267, 1, 
/* out0247_had-eta7-phi12*/	4, 61, 1, 62, 5, 75, 1, 266, 3, 
/* out0248_had-eta8-phi12*/	6, 61, 4, 75, 2, 174, 5, 180, 2, 234, 3, 266, 2, 
/* out0249_had-eta9-phi12*/	7, 61, 1, 74, 3, 173, 4, 174, 2, 180, 2, 234, 6, 266, 1, 
/* out0250_had-eta10-phi12*/	5, 60, 1, 74, 3, 173, 5, 233, 4, 234, 2, 
/* out0251_had-eta11-phi12*/	3, 20, 3, 172, 4, 233, 4, 
/* out0252_had-eta12-phi12*/	5, 20, 3, 172, 4, 228, 2, 232, 1, 233, 1, 
/* out0253_had-eta13-phi12*/	6, 19, 2, 20, 1, 171, 2, 172, 1, 228, 1, 232, 2, 
/* out0254_had-eta14-phi12*/	3, 19, 2, 171, 2, 227, 2, 
/* out0255_had-eta15-phi12*/	4, 19, 2, 166, 1, 171, 1, 227, 2, 
/* out0256_had-eta16-phi12*/	6, 18, 1, 19, 1, 166, 1, 170, 1, 226, 2, 227, 1, 
/* out0257_had-eta17-phi12*/	3, 18, 1, 170, 1, 226, 3, 
/* out0258_had-eta18-phi12*/	1, 18, 1, 
/* out0259_had-eta19-phi12*/	2, 4, 1, 18, 1, 
/* out0260_had-eta0-phi13*/	1, 273, 1, 
/* out0261_had-eta1-phi13*/	1, 273, 5, 
/* out0262_had-eta2-phi13*/	5, 65, 1, 66, 11, 79, 4, 272, 2, 273, 2, 
/* out0263_had-eta3-phi13*/	4, 65, 7, 78, 4, 79, 3, 272, 4, 
/* out0264_had-eta4-phi13*/	5, 64, 5, 77, 3, 78, 4, 271, 3, 272, 2, 
/* out0265_had-eta5-phi13*/	4, 63, 2, 76, 1, 77, 7, 271, 4, 
/* out0266_had-eta6-phi13*/	3, 76, 8, 270, 2, 271, 1, 
/* out0267_had-eta7-phi13*/	3, 75, 5, 76, 2, 270, 3, 
/* out0268_had-eta8-phi13*/	5, 75, 6, 174, 6, 230, 3, 234, 1, 270, 2, 
/* out0269_had-eta9-phi13*/	8, 74, 5, 169, 3, 173, 3, 174, 3, 229, 2, 230, 5, 234, 2, 270, 1, 
/* out0270_had-eta10-phi13*/	4, 74, 4, 168, 1, 173, 4, 229, 5, 
/* out0271_had-eta11-phi13*/	5, 20, 3, 168, 3, 172, 1, 228, 2, 229, 2, 
/* out0272_had-eta12-phi13*/	5, 20, 3, 167, 1, 168, 1, 172, 2, 228, 4, 
/* out0273_had-eta13-phi13*/	6, 7, 1, 19, 1, 20, 1, 167, 3, 227, 1, 228, 2, 
/* out0274_had-eta14-phi13*/	4, 19, 1, 167, 2, 171, 1, 227, 3, 
/* out0275_had-eta15-phi13*/	4, 6, 1, 19, 1, 166, 2, 227, 2, 
/* out0276_had-eta16-phi13*/	4, 6, 1, 166, 2, 226, 2, 227, 1, 
/* out0277_had-eta17-phi13*/	3, 6, 1, 166, 1, 226, 3, 
/* out0278_had-eta18-phi13*/	3, 4, 1, 18, 1, 226, 1, 
/* out0279_had-eta19-phi13*/	1, 4, 2, 
/* out0280_had-eta0-phi14*/	1, 273, 1, 
/* out0281_had-eta1-phi14*/	1, 273, 5, 
/* out0282_had-eta2-phi14*/	3, 79, 5, 272, 2, 273, 2, 
/* out0283_had-eta3-phi14*/	3, 78, 4, 79, 4, 272, 4, 
/* out0284_had-eta4-phi14*/	5, 33, 7, 77, 2, 78, 4, 271, 3, 272, 2, 
/* out0285_had-eta5-phi14*/	4, 32, 5, 33, 1, 77, 4, 271, 4, 
/* out0286_had-eta6-phi14*/	5, 31, 2, 32, 3, 76, 3, 270, 2, 271, 1, 
/* out0287_had-eta7-phi14*/	4, 31, 5, 75, 1, 76, 1, 270, 3, 
/* out0288_had-eta8-phi14*/	5, 30, 4, 75, 1, 169, 3, 230, 2, 270, 2, 
/* out0289_had-eta9-phi14*/	7, 30, 4, 74, 1, 169, 6, 225, 2, 229, 1, 230, 6, 270, 1, 
/* out0290_had-eta10-phi14*/	5, 29, 4, 168, 3, 169, 2, 225, 1, 229, 5, 
/* out0291_had-eta11-phi14*/	5, 29, 3, 168, 4, 224, 2, 228, 1, 229, 1, 
/* out0292_had-eta12-phi14*/	5, 7, 2, 29, 1, 167, 2, 168, 1, 228, 3, 
/* out0293_had-eta13-phi14*/	4, 7, 2, 167, 3, 223, 2, 228, 1, 
/* out0294_had-eta14-phi14*/	4, 7, 2, 167, 2, 223, 1, 227, 2, 
/* out0295_had-eta15-phi14*/	3, 6, 2, 166, 2, 227, 2, 
/* out0296_had-eta16-phi14*/	3, 6, 1, 166, 2, 222, 1, 
/* out0297_had-eta17-phi14*/	4, 6, 1, 166, 2, 222, 1, 226, 2, 
/* out0298_had-eta18-phi14*/	3, 4, 1, 6, 1, 226, 1, 
/* out0299_had-eta19-phi14*/	1, 4, 3, 
/* out0300_had-eta0-phi15*/	1, 277, 1, 
/* out0301_had-eta1-phi15*/	1, 277, 5, 
/* out0302_had-eta2-phi15*/	3, 45, 5, 276, 2, 277, 2, 
/* out0303_had-eta3-phi15*/	3, 44, 4, 45, 4, 276, 4, 
/* out0304_had-eta4-phi15*/	5, 33, 7, 43, 2, 44, 4, 275, 3, 276, 2, 
/* out0305_had-eta5-phi15*/	4, 32, 5, 33, 1, 43, 4, 275, 4, 
/* out0306_had-eta6-phi15*/	5, 31, 2, 32, 3, 42, 3, 274, 2, 275, 1, 
/* out0307_had-eta7-phi15*/	4, 31, 6, 41, 1, 42, 1, 274, 3, 
/* out0308_had-eta8-phi15*/	6, 30, 4, 31, 1, 41, 1, 165, 5, 225, 1, 274, 2, 
/* out0309_had-eta9-phi15*/	7, 30, 4, 40, 1, 164, 2, 165, 3, 169, 2, 225, 6, 274, 1, 
/* out0310_had-eta10-phi15*/	5, 29, 4, 164, 4, 168, 1, 224, 2, 225, 3, 
/* out0311_had-eta11-phi15*/	5, 29, 3, 163, 2, 164, 1, 168, 2, 224, 5, 
/* out0312_had-eta12-phi15*/	5, 7, 2, 29, 1, 163, 3, 223, 1, 224, 2, 
/* out0313_had-eta13-phi15*/	5, 7, 3, 162, 1, 163, 1, 167, 2, 223, 3, 
/* out0314_had-eta14-phi15*/	4, 7, 2, 162, 2, 167, 1, 223, 3, 
/* out0315_had-eta15-phi15*/	4, 6, 2, 162, 1, 166, 1, 222, 2, 
/* out0316_had-eta16-phi15*/	3, 6, 1, 166, 1, 222, 2, 
/* out0317_had-eta17-phi15*/	4, 6, 1, 161, 2, 166, 1, 222, 2, 
/* out0318_had-eta18-phi15*/	2, 4, 1, 6, 1, 
/* out0319_had-eta19-phi15*/	1, 4, 3, 
/* out0320_had-eta0-phi16*/	1, 277, 1, 
/* out0321_had-eta1-phi16*/	1, 277, 5, 
/* out0322_had-eta2-phi16*/	5, 45, 4, 58, 1, 59, 11, 276, 2, 277, 2, 
/* out0323_had-eta3-phi16*/	4, 44, 4, 45, 3, 58, 7, 276, 4, 
/* out0324_had-eta4-phi16*/	5, 43, 3, 44, 4, 57, 5, 275, 3, 276, 2, 
/* out0325_had-eta5-phi16*/	4, 42, 1, 43, 7, 56, 2, 275, 4, 
/* out0326_had-eta6-phi16*/	3, 42, 8, 274, 2, 275, 1, 
/* out0327_had-eta7-phi16*/	3, 41, 5, 42, 2, 274, 3, 
/* out0328_had-eta8-phi16*/	5, 41, 6, 160, 1, 165, 5, 221, 4, 274, 2, 
/* out0329_had-eta9-phi16*/	8, 40, 5, 160, 2, 164, 3, 165, 3, 220, 2, 221, 5, 225, 2, 274, 1, 
/* out0330_had-eta10-phi16*/	5, 40, 4, 164, 5, 220, 4, 224, 1, 225, 1, 
/* out0331_had-eta11-phi16*/	6, 13, 3, 163, 3, 164, 1, 219, 1, 220, 1, 224, 3, 
/* out0332_had-eta12-phi16*/	5, 13, 3, 163, 3, 219, 2, 223, 1, 224, 1, 
/* out0333_had-eta13-phi16*/	6, 7, 1, 11, 1, 13, 1, 162, 2, 163, 1, 223, 3, 
/* out0334_had-eta14-phi16*/	4, 7, 1, 11, 1, 162, 2, 223, 2, 
/* out0335_had-eta15-phi16*/	4, 6, 1, 11, 1, 162, 2, 222, 2, 
/* out0336_had-eta16-phi16*/	4, 6, 1, 161, 2, 162, 1, 222, 2, 
/* out0337_had-eta17-phi16*/	3, 6, 1, 161, 3, 222, 2, 
/* out0338_had-eta18-phi16*/	2, 4, 1, 5, 1, 
/* out0339_had-eta19-phi16*/	1, 4, 2, 
/* out0340_had-eta0-phi17*/	1, 281, 1, 
/* out0341_had-eta1-phi17*/	1, 281, 5, 
/* out0342_had-eta2-phi17*/	5, 58, 1, 59, 5, 97, 10, 280, 2, 281, 2, 
/* out0343_had-eta3-phi17*/	5, 57, 1, 58, 7, 96, 6, 97, 2, 280, 4, 
/* out0344_had-eta4-phi17*/	5, 57, 10, 95, 2, 96, 1, 279, 3, 280, 2, 
/* out0345_had-eta5-phi17*/	3, 56, 10, 95, 1, 279, 4, 
/* out0346_had-eta6-phi17*/	5, 42, 1, 55, 5, 56, 3, 278, 2, 279, 1, 
/* out0347_had-eta7-phi17*/	4, 41, 1, 54, 1, 55, 5, 278, 3, 
/* out0348_had-eta8-phi17*/	6, 41, 2, 54, 4, 160, 4, 216, 1, 221, 4, 278, 2, 
/* out0349_had-eta9-phi17*/	7, 40, 3, 54, 1, 160, 6, 216, 2, 220, 3, 221, 3, 278, 1, 
/* out0350_had-eta10-phi17*/	4, 40, 3, 53, 1, 158, 5, 220, 5, 
/* out0351_had-eta11-phi17*/	5, 13, 3, 158, 4, 163, 1, 219, 3, 220, 1, 
/* out0352_had-eta12-phi17*/	4, 13, 3, 156, 2, 163, 2, 219, 4, 
/* out0353_had-eta13-phi17*/	6, 11, 2, 13, 1, 156, 2, 162, 1, 218, 1, 219, 1, 
/* out0354_had-eta14-phi17*/	3, 11, 2, 162, 2, 218, 3, 
/* out0355_had-eta15-phi17*/	3, 11, 2, 162, 2, 218, 2, 
/* out0356_had-eta16-phi17*/	5, 5, 1, 11, 1, 161, 3, 217, 1, 222, 1, 
/* out0357_had-eta17-phi17*/	4, 5, 1, 161, 3, 217, 1, 222, 1, 
/* out0358_had-eta18-phi17*/	1, 5, 1, 
/* out0359_had-eta19-phi17*/	2, 4, 1, 5, 1, 
/* out0360_had-eta0-phi18*/	1, 281, 1, 
/* out0361_had-eta1-phi18*/	1, 281, 5, 
/* out0362_had-eta2-phi18*/	5, 97, 4, 110, 7, 111, 1, 280, 2, 281, 2, 
/* out0363_had-eta3-phi18*/	4, 96, 7, 108, 3, 110, 4, 280, 4, 
/* out0364_had-eta4-phi18*/	5, 95, 9, 96, 2, 108, 2, 279, 3, 280, 2, 
/* out0365_had-eta5-phi18*/	4, 56, 1, 94, 5, 95, 4, 279, 4, 
/* out0366_had-eta6-phi18*/	5, 55, 3, 93, 1, 94, 5, 278, 2, 279, 1, 
/* out0367_had-eta7-phi18*/	4, 54, 1, 55, 3, 93, 3, 278, 3, 
/* out0368_had-eta8-phi18*/	5, 54, 6, 159, 1, 160, 1, 216, 3, 278, 2, 
/* out0369_had-eta9-phi18*/	6, 53, 2, 54, 2, 159, 4, 160, 2, 216, 7, 278, 1, 
/* out0370_had-eta10-phi18*/	4, 53, 4, 158, 4, 159, 1, 214, 5, 
/* out0371_had-eta11-phi18*/	5, 13, 1, 53, 2, 158, 3, 214, 3, 219, 1, 
/* out0372_had-eta12-phi18*/	5, 12, 2, 13, 1, 156, 4, 213, 1, 219, 3, 
/* out0373_had-eta13-phi18*/	6, 11, 1, 12, 1, 156, 3, 213, 1, 218, 2, 219, 1, 
/* out0374_had-eta14-phi18*/	4, 11, 2, 155, 2, 156, 1, 218, 3, 
/* out0375_had-eta15-phi18*/	3, 11, 2, 155, 2, 218, 2, 
/* out0376_had-eta16-phi18*/	4, 5, 1, 155, 1, 161, 1, 217, 2, 
/* out0377_had-eta17-phi18*/	3, 5, 1, 161, 2, 217, 2, 
/* out0378_had-eta18-phi18*/	2, 5, 1, 217, 1, 
/* out0379_had-eta19-phi18*/	1, 5, 1, 
/* out0380_had-eta0-phi19*/	1, 285, 1, 
/* out0381_had-eta1-phi19*/	1, 285, 5, 
/* out0382_had-eta2-phi19*/	5, 109, 4, 110, 3, 111, 15, 284, 2, 285, 2, 
/* out0383_had-eta3-phi19*/	5, 107, 1, 108, 7, 109, 6, 110, 2, 284, 4, 
/* out0384_had-eta4-phi19*/	5, 106, 7, 107, 1, 108, 4, 283, 3, 284, 2, 
/* out0385_had-eta5-phi19*/	4, 94, 3, 105, 2, 106, 6, 283, 4, 
/* out0386_had-eta6-phi19*/	5, 93, 3, 94, 3, 105, 3, 282, 2, 283, 1, 
/* out0387_had-eta7-phi19*/	2, 93, 7, 282, 3, 
/* out0388_had-eta8-phi19*/	7, 54, 1, 92, 4, 93, 1, 159, 1, 215, 1, 216, 1, 282, 2, 
/* out0389_had-eta9-phi19*/	6, 53, 2, 92, 3, 159, 6, 215, 6, 216, 2, 282, 1, 
/* out0390_had-eta10-phi19*/	5, 53, 4, 157, 3, 159, 2, 214, 5, 215, 1, 
/* out0391_had-eta11-phi19*/	5, 12, 2, 53, 1, 157, 4, 213, 1, 214, 3, 
/* out0392_had-eta12-phi19*/	4, 12, 3, 156, 2, 157, 1, 213, 4, 
/* out0393_had-eta13-phi19*/	4, 12, 2, 156, 2, 194, 1, 213, 3, 
/* out0394_had-eta14-phi19*/	5, 11, 1, 16, 1, 155, 3, 207, 1, 218, 2, 
/* out0395_had-eta15-phi19*/	4, 16, 1, 155, 2, 207, 1, 218, 1, 
/* out0396_had-eta16-phi19*/	3, 5, 1, 155, 2, 217, 2, 
/* out0397_had-eta17-phi19*/	2, 5, 1, 217, 2, 
/* out0398_had-eta18-phi19*/	2, 5, 1, 217, 1, 
/* out0399_had-eta19-phi19*/	1, 5, 1, 
/* out0400_had-eta0-phi20*/	1, 285, 1, 
/* out0401_had-eta1-phi20*/	1, 285, 5, 
/* out0402_had-eta2-phi20*/	4, 109, 3, 121, 2, 284, 2, 285, 2, 
/* out0403_had-eta3-phi20*/	4, 107, 7, 109, 3, 121, 6, 284, 4, 
/* out0404_had-eta4-phi20*/	5, 106, 2, 107, 7, 117, 4, 283, 3, 284, 2, 
/* out0405_had-eta5-phi20*/	4, 105, 4, 106, 1, 117, 4, 283, 4, 
/* out0406_had-eta6-phi20*/	4, 105, 7, 127, 1, 282, 2, 283, 1, 
/* out0407_had-eta7-phi20*/	3, 93, 1, 127, 6, 282, 3, 
/* out0408_had-eta8-phi20*/	3, 92, 5, 127, 1, 282, 2, 
/* out0409_had-eta9-phi20*/	6, 92, 4, 132, 1, 159, 1, 197, 5, 215, 7, 282, 1, 
/* out0410_had-eta10-phi20*/	5, 132, 4, 157, 3, 197, 2, 211, 4, 215, 1, 
/* out0411_had-eta11-phi20*/	5, 12, 1, 132, 2, 157, 4, 211, 4, 213, 1, 
/* out0412_had-eta12-phi20*/	4, 12, 3, 157, 1, 194, 3, 213, 3, 
/* out0413_had-eta13-phi20*/	5, 12, 2, 16, 1, 194, 3, 207, 1, 213, 2, 
/* out0414_had-eta14-phi20*/	4, 16, 2, 155, 1, 194, 1, 207, 2, 
/* out0415_had-eta15-phi20*/	3, 16, 2, 155, 2, 207, 2, 
/* out0416_had-eta16-phi20*/	4, 16, 1, 155, 1, 207, 1, 217, 1, 
/* out0417_had-eta17-phi20*/	2, 5, 1, 217, 2, 
/* out0418_had-eta18-phi20*/	2, 5, 1, 217, 1, 
/* out0419_had-eta19-phi20*/	1, 5, 1, 
/* out0420_had-eta0-phi21*/	1, 289, 1, 
/* out0421_had-eta1-phi21*/	1, 289, 5, 
/* out0422_had-eta2-phi21*/	4, 119, 3, 121, 2, 288, 2, 289, 2, 
/* out0423_had-eta3-phi21*/	4, 118, 7, 119, 3, 121, 6, 288, 4, 
/* out0424_had-eta4-phi21*/	5, 117, 4, 118, 7, 129, 2, 287, 3, 288, 2, 
/* out0425_had-eta5-phi21*/	4, 117, 4, 128, 4, 129, 1, 287, 4, 
/* out0426_had-eta6-phi21*/	4, 127, 1, 128, 7, 286, 2, 287, 1, 
/* out0427_had-eta7-phi21*/	3, 127, 6, 134, 1, 286, 3, 
/* out0428_had-eta8-phi21*/	4, 127, 1, 133, 5, 197, 1, 286, 2, 
/* out0429_had-eta9-phi21*/	6, 132, 1, 133, 4, 196, 1, 197, 5, 212, 7, 286, 1, 
/* out0430_had-eta10-phi21*/	5, 132, 4, 195, 3, 197, 3, 211, 4, 212, 1, 
/* out0431_had-eta11-phi21*/	5, 17, 1, 132, 3, 195, 4, 208, 1, 211, 4, 
/* out0432_had-eta12-phi21*/	4, 17, 3, 194, 3, 195, 1, 208, 3, 
/* out0433_had-eta13-phi21*/	5, 16, 1, 17, 2, 194, 3, 207, 1, 208, 2, 
/* out0434_had-eta14-phi21*/	4, 16, 2, 151, 1, 194, 1, 207, 2, 
/* out0435_had-eta15-phi21*/	3, 16, 2, 151, 2, 207, 2, 
/* out0436_had-eta16-phi21*/	4, 16, 1, 151, 1, 202, 1, 207, 1, 
/* out0437_had-eta17-phi21*/	2, 21, 1, 202, 2, 
/* out0438_had-eta18-phi21*/	2, 21, 1, 202, 1, 
/* out0439_had-eta19-phi21*/	1, 21, 1, 
/* out0440_had-eta0-phi22*/	1, 289, 1, 
/* out0441_had-eta1-phi22*/	1, 289, 5, 
/* out0442_had-eta2-phi22*/	5, 119, 4, 120, 15, 131, 3, 288, 2, 289, 2, 
/* out0443_had-eta3-phi22*/	5, 118, 1, 119, 6, 130, 7, 131, 2, 288, 4, 
/* out0444_had-eta4-phi22*/	5, 118, 1, 129, 7, 130, 4, 287, 3, 288, 2, 
/* out0445_had-eta5-phi22*/	4, 128, 2, 129, 6, 135, 3, 287, 4, 
/* out0446_had-eta6-phi22*/	5, 128, 3, 134, 3, 135, 3, 286, 2, 287, 1, 
/* out0447_had-eta7-phi22*/	2, 134, 7, 286, 3, 
/* out0448_had-eta8-phi22*/	7, 68, 1, 133, 4, 134, 1, 196, 1, 210, 1, 212, 1, 286, 2, 
/* out0449_had-eta9-phi22*/	6, 67, 2, 133, 3, 196, 6, 210, 2, 212, 6, 286, 1, 
/* out0450_had-eta10-phi22*/	6, 67, 4, 132, 1, 195, 3, 196, 2, 209, 5, 212, 1, 
/* out0451_had-eta11-phi22*/	5, 17, 2, 67, 1, 195, 4, 208, 1, 209, 3, 
/* out0452_had-eta12-phi22*/	4, 17, 3, 152, 2, 195, 1, 208, 4, 
/* out0453_had-eta13-phi22*/	4, 17, 2, 152, 2, 194, 1, 208, 3, 
/* out0454_had-eta14-phi22*/	5, 16, 1, 22, 1, 151, 3, 203, 2, 207, 1, 
/* out0455_had-eta15-phi22*/	4, 16, 1, 151, 2, 203, 1, 207, 1, 
/* out0456_had-eta16-phi22*/	3, 21, 1, 151, 2, 202, 2, 
/* out0457_had-eta17-phi22*/	2, 21, 1, 202, 2, 
/* out0458_had-eta18-phi22*/	2, 21, 1, 202, 1, 
/* out0459_had-eta19-phi22*/	1, 21, 1, 
/* out0460_had-eta0-phi23*/	1, 293, 1, 
/* out0461_had-eta1-phi23*/	1, 293, 5, 
/* out0462_had-eta2-phi23*/	5, 120, 1, 131, 7, 138, 4, 292, 2, 293, 2, 
/* out0463_had-eta3-phi23*/	4, 130, 3, 131, 4, 137, 7, 292, 4, 
/* out0464_had-eta4-phi23*/	5, 130, 2, 136, 9, 137, 2, 291, 3, 292, 2, 
/* out0465_had-eta5-phi23*/	4, 70, 1, 135, 5, 136, 4, 291, 4, 
/* out0466_had-eta6-phi23*/	5, 69, 3, 134, 1, 135, 5, 290, 2, 291, 1, 
/* out0467_had-eta7-phi23*/	4, 68, 1, 69, 3, 134, 3, 290, 3, 
/* out0468_had-eta8-phi23*/	5, 68, 6, 154, 1, 196, 1, 210, 3, 290, 2, 
/* out0469_had-eta9-phi23*/	6, 67, 2, 68, 2, 154, 2, 196, 4, 210, 7, 290, 1, 
/* out0470_had-eta10-phi23*/	4, 67, 4, 153, 4, 196, 1, 209, 5, 
/* out0471_had-eta11-phi23*/	5, 23, 1, 67, 2, 153, 3, 204, 1, 209, 3, 
/* out0472_had-eta12-phi23*/	5, 17, 2, 23, 1, 152, 4, 204, 3, 208, 1, 
/* out0473_had-eta13-phi23*/	6, 17, 1, 22, 1, 152, 3, 203, 2, 204, 1, 208, 1, 
/* out0474_had-eta14-phi23*/	4, 22, 2, 151, 2, 152, 1, 203, 3, 
/* out0475_had-eta15-phi23*/	3, 22, 2, 151, 2, 203, 2, 
/* out0476_had-eta16-phi23*/	4, 21, 1, 146, 1, 151, 1, 202, 2, 
/* out0477_had-eta17-phi23*/	3, 21, 1, 146, 2, 202, 2, 
/* out0478_had-eta18-phi23*/	2, 21, 1, 202, 1, 
/* out0479_had-eta19-phi23*/	1, 21, 1, 
/* out0480_had-eta0-phi24*/	1, 293, 1, 
/* out0481_had-eta1-phi24*/	1, 293, 5, 
/* out0482_had-eta2-phi24*/	5, 72, 1, 73, 5, 138, 10, 292, 2, 293, 2, 
/* out0483_had-eta3-phi24*/	5, 71, 1, 72, 7, 137, 6, 138, 2, 292, 4, 
/* out0484_had-eta4-phi24*/	5, 71, 10, 136, 2, 137, 1, 291, 3, 292, 2, 
/* out0485_had-eta5-phi24*/	3, 70, 10, 136, 1, 291, 4, 
/* out0486_had-eta6-phi24*/	5, 69, 5, 70, 3, 82, 1, 290, 2, 291, 1, 
/* out0487_had-eta7-phi24*/	4, 68, 1, 69, 5, 81, 1, 290, 3, 
/* out0488_had-eta8-phi24*/	6, 68, 4, 81, 2, 154, 4, 206, 4, 210, 1, 290, 2, 
/* out0489_had-eta9-phi24*/	7, 68, 1, 80, 3, 154, 6, 205, 3, 206, 3, 210, 2, 290, 1, 
/* out0490_had-eta10-phi24*/	4, 67, 1, 80, 3, 153, 5, 205, 5, 
/* out0491_had-eta11-phi24*/	5, 23, 3, 148, 1, 153, 4, 204, 3, 205, 1, 
/* out0492_had-eta12-phi24*/	4, 23, 3, 148, 2, 152, 2, 204, 4, 
/* out0493_had-eta13-phi24*/	6, 22, 2, 23, 1, 147, 1, 152, 2, 203, 1, 204, 1, 
/* out0494_had-eta14-phi24*/	3, 22, 2, 147, 2, 203, 3, 
/* out0495_had-eta15-phi24*/	3, 22, 2, 147, 2, 203, 2, 
/* out0496_had-eta16-phi24*/	5, 21, 1, 22, 1, 146, 3, 198, 1, 202, 1, 
/* out0497_had-eta17-phi24*/	4, 21, 1, 146, 3, 198, 1, 202, 1, 
/* out0498_had-eta18-phi24*/	1, 21, 1, 
/* out0499_had-eta19-phi24*/	1, 21, 1, 
/* out0500_had-eta0-phi25*/	1, 297, 1, 
/* out0501_had-eta1-phi25*/	1, 297, 5, 
/* out0502_had-eta2-phi25*/	5, 72, 1, 73, 11, 85, 4, 296, 2, 297, 2, 
/* out0503_had-eta3-phi25*/	4, 72, 7, 84, 4, 85, 3, 296, 4, 
/* out0504_had-eta4-phi25*/	5, 71, 5, 83, 3, 84, 4, 295, 3, 296, 2, 
/* out0505_had-eta5-phi25*/	4, 70, 2, 82, 1, 83, 7, 295, 4, 
/* out0506_had-eta6-phi25*/	3, 82, 8, 294, 2, 295, 1, 
/* out0507_had-eta7-phi25*/	3, 81, 5, 82, 2, 294, 3, 
/* out0508_had-eta8-phi25*/	5, 81, 6, 150, 5, 154, 1, 206, 4, 294, 2, 
/* out0509_had-eta9-phi25*/	8, 80, 5, 149, 3, 150, 3, 154, 2, 201, 2, 205, 2, 206, 5, 294, 1, 
/* out0510_had-eta10-phi25*/	5, 80, 4, 149, 5, 200, 1, 201, 1, 205, 4, 
/* out0511_had-eta11-phi25*/	6, 23, 3, 148, 3, 149, 1, 200, 3, 204, 1, 205, 1, 
/* out0512_had-eta12-phi25*/	5, 23, 3, 148, 3, 199, 1, 200, 1, 204, 2, 
/* out0513_had-eta13-phi25*/	5, 22, 1, 23, 1, 147, 2, 148, 1, 199, 3, 
/* out0514_had-eta14-phi25*/	3, 22, 1, 147, 2, 199, 2, 
/* out0515_had-eta15-phi25*/	3, 22, 1, 147, 2, 198, 2, 
/* out0516_had-eta16-phi25*/	3, 146, 2, 147, 1, 198, 2, 
/* out0517_had-eta17-phi25*/	2, 146, 3, 198, 2, 
/* out0518_had-eta18-phi25*/	1, 21, 1, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	1, 297, 1, 
/* out0521_had-eta1-phi26*/	1, 297, 5, 
/* out0522_had-eta2-phi26*/	3, 85, 5, 296, 2, 297, 2, 
/* out0523_had-eta3-phi26*/	3, 84, 4, 85, 4, 296, 4, 
/* out0524_had-eta4-phi26*/	4, 83, 2, 84, 4, 295, 3, 296, 2, 
/* out0525_had-eta5-phi26*/	2, 83, 4, 295, 4, 
/* out0526_had-eta6-phi26*/	3, 82, 3, 294, 2, 295, 1, 
/* out0527_had-eta7-phi26*/	3, 81, 1, 82, 1, 294, 3, 
/* out0528_had-eta8-phi26*/	4, 81, 1, 150, 5, 201, 1, 294, 2, 
/* out0529_had-eta9-phi26*/	5, 80, 1, 149, 2, 150, 3, 201, 6, 294, 1, 
/* out0530_had-eta10-phi26*/	3, 149, 4, 200, 2, 201, 3, 
/* out0531_had-eta11-phi26*/	3, 148, 2, 149, 1, 200, 5, 
/* out0532_had-eta12-phi26*/	3, 148, 3, 199, 1, 200, 2, 
/* out0533_had-eta13-phi26*/	3, 147, 1, 148, 1, 199, 3, 
/* out0534_had-eta14-phi26*/	2, 147, 2, 199, 3, 
/* out0535_had-eta15-phi26*/	2, 147, 1, 198, 2, 
/* out0536_had-eta16-phi26*/	1, 198, 2, 
/* out0537_had-eta17-phi26*/	2, 146, 2, 198, 2, 
/* out0538_had-eta18-phi26*/	0, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	1, 201, 2, 
/* out0550_had-eta10-phi27*/	1, 201, 1, 
/* out0551_had-eta11-phi27*/	1, 200, 2, 
/* out0552_had-eta12-phi27*/	0, 
/* out0553_had-eta13-phi27*/	1, 199, 2, 
/* out0554_had-eta14-phi27*/	1, 199, 1, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	1, 198, 1, 
/* out0557_had-eta17-phi27*/	1, 198, 1, 
/* out0558_had-eta18-phi27*/	0, 
/* out0559_had-eta19-phi27*/	0, 
};