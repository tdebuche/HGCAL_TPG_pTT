parameter integer matrixH [0:2618] = {
/* num inputs = 180(in0-in179) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 4 */
//* total number of input in adders 1069 */

/* out0000_had-eta0-phi0*/	1, 135, 3, 
/* out0001_had-eta1-phi0*/	1, 135, 4, 
/* out0002_had-eta2-phi0*/	2, 134, 4, 135, 1, 
/* out0003_had-eta3-phi0*/	1, 134, 4, 
/* out0004_had-eta4-phi0*/	1, 133, 4, 
/* out0005_had-eta5-phi0*/	3, 87, 11, 94, 1, 133, 4, 
/* out0006_had-eta6-phi0*/	3, 86, 6, 87, 4, 132, 3, 
/* out0007_had-eta7-phi0*/	3, 85, 1, 86, 8, 132, 3, 
/* out0008_had-eta8-phi0*/	2, 85, 8, 132, 2, 
/* out0009_had-eta9-phi0*/	2, 84, 3, 85, 3, 
/* out0010_had-eta10-phi0*/	1, 84, 5, 
/* out0011_had-eta11-phi0*/	3, 83, 2, 84, 3, 127, 3, 
/* out0012_had-eta12-phi0*/	3, 83, 4, 126, 1, 127, 4, 
/* out0013_had-eta13-phi0*/	2, 83, 3, 126, 3, 
/* out0014_had-eta14-phi0*/	2, 82, 2, 126, 1, 
/* out0015_had-eta15-phi0*/	2, 82, 2, 125, 2, 
/* out0016_had-eta16-phi0*/	2, 82, 2, 125, 2, 
/* out0017_had-eta17-phi0*/	2, 81, 2, 82, 1, 
/* out0018_had-eta18-phi0*/	2, 81, 3, 124, 2, 
/* out0019_had-eta19-phi0*/	2, 81, 1, 124, 1, 
/* out0020_had-eta0-phi1*/	1, 135, 3, 
/* out0021_had-eta1-phi1*/	1, 135, 4, 
/* out0022_had-eta2-phi1*/	2, 134, 4, 135, 1, 
/* out0023_had-eta3-phi1*/	1, 134, 4, 
/* out0024_had-eta4-phi1*/	1, 133, 4, 
/* out0025_had-eta5-phi1*/	4, 87, 1, 93, 3, 94, 14, 133, 4, 
/* out0026_had-eta6-phi1*/	3, 86, 1, 93, 9, 132, 3, 
/* out0027_had-eta7-phi1*/	3, 86, 1, 92, 7, 132, 3, 
/* out0028_had-eta8-phi1*/	4, 85, 3, 91, 1, 92, 2, 132, 2, 
/* out0029_had-eta9-phi1*/	3, 84, 1, 85, 1, 91, 4, 
/* out0030_had-eta10-phi1*/	3, 84, 3, 90, 1, 91, 1, 
/* out0031_had-eta11-phi1*/	4, 83, 1, 84, 1, 90, 2, 127, 4, 
/* out0032_had-eta12-phi1*/	3, 83, 3, 126, 2, 127, 5, 
/* out0033_had-eta13-phi1*/	2, 83, 3, 126, 4, 
/* out0034_had-eta14-phi1*/	3, 82, 2, 125, 1, 126, 2, 
/* out0035_had-eta15-phi1*/	2, 82, 2, 125, 3, 
/* out0036_had-eta16-phi1*/	2, 82, 2, 125, 2, 
/* out0037_had-eta17-phi1*/	3, 81, 2, 124, 1, 125, 1, 
/* out0038_had-eta18-phi1*/	2, 81, 2, 124, 3, 
/* out0039_had-eta19-phi1*/	2, 81, 1, 124, 1, 
/* out0040_had-eta0-phi2*/	1, 139, 3, 
/* out0041_had-eta1-phi2*/	1, 139, 4, 
/* out0042_had-eta2-phi2*/	2, 138, 4, 139, 1, 
/* out0043_had-eta3-phi2*/	1, 138, 4, 
/* out0044_had-eta4-phi2*/	1, 137, 4, 
/* out0045_had-eta5-phi2*/	4, 70, 12, 93, 1, 94, 1, 137, 4, 
/* out0046_had-eta6-phi2*/	4, 69, 6, 70, 1, 93, 3, 136, 3, 
/* out0047_had-eta7-phi2*/	4, 68, 1, 69, 2, 92, 5, 136, 3, 
/* out0048_had-eta8-phi2*/	4, 68, 2, 91, 3, 92, 2, 136, 2, 
/* out0049_had-eta9-phi2*/	1, 91, 5, 
/* out0050_had-eta10-phi2*/	2, 90, 3, 91, 1, 
/* out0051_had-eta11-phi2*/	2, 90, 4, 122, 3, 
/* out0052_had-eta12-phi2*/	3, 89, 1, 90, 1, 122, 4, 
/* out0053_had-eta13-phi2*/	4, 89, 3, 121, 1, 122, 1, 126, 2, 
/* out0054_had-eta14-phi2*/	3, 89, 2, 121, 2, 126, 1, 
/* out0055_had-eta15-phi2*/	3, 82, 2, 121, 1, 125, 2, 
/* out0056_had-eta16-phi2*/	3, 82, 1, 88, 1, 125, 2, 
/* out0057_had-eta17-phi2*/	4, 81, 2, 88, 1, 124, 2, 125, 1, 
/* out0058_had-eta18-phi2*/	2, 81, 2, 124, 3, 
/* out0059_had-eta19-phi2*/	1, 124, 1, 
/* out0060_had-eta0-phi3*/	1, 139, 3, 
/* out0061_had-eta1-phi3*/	1, 139, 4, 
/* out0062_had-eta2-phi3*/	2, 138, 4, 139, 1, 
/* out0063_had-eta3-phi3*/	1, 138, 4, 
/* out0064_had-eta4-phi3*/	1, 137, 4, 
/* out0065_had-eta5-phi3*/	3, 70, 3, 73, 6, 137, 4, 
/* out0066_had-eta6-phi3*/	4, 69, 6, 72, 1, 73, 2, 136, 3, 
/* out0067_had-eta7-phi3*/	4, 68, 4, 69, 2, 72, 1, 136, 3, 
/* out0068_had-eta8-phi3*/	2, 68, 6, 136, 2, 
/* out0069_had-eta9-phi3*/	2, 67, 5, 91, 1, 
/* out0070_had-eta10-phi3*/	2, 67, 3, 90, 1, 
/* out0071_had-eta11-phi3*/	3, 66, 1, 90, 3, 122, 3, 
/* out0072_had-eta12-phi3*/	4, 66, 1, 89, 2, 90, 1, 122, 4, 
/* out0073_had-eta13-phi3*/	3, 89, 3, 121, 3, 122, 1, 
/* out0074_had-eta14-phi3*/	2, 89, 2, 121, 3, 
/* out0075_had-eta15-phi3*/	3, 88, 2, 120, 1, 121, 2, 
/* out0076_had-eta16-phi3*/	2, 88, 2, 120, 2, 
/* out0077_had-eta17-phi3*/	2, 88, 1, 120, 2, 
/* out0078_had-eta18-phi3*/	2, 81, 1, 124, 2, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	1, 143, 3, 
/* out0081_had-eta1-phi4*/	1, 143, 4, 
/* out0082_had-eta2-phi4*/	2, 142, 4, 143, 1, 
/* out0083_had-eta3-phi4*/	1, 142, 4, 
/* out0084_had-eta4-phi4*/	1, 141, 4, 
/* out0085_had-eta5-phi4*/	3, 73, 6, 74, 2, 141, 4, 
/* out0086_had-eta6-phi4*/	4, 72, 6, 73, 2, 74, 2, 140, 3, 
/* out0087_had-eta7-phi4*/	4, 68, 1, 71, 1, 72, 6, 140, 3, 
/* out0088_had-eta8-phi4*/	3, 68, 2, 71, 5, 140, 2, 
/* out0089_had-eta9-phi4*/	2, 67, 5, 71, 1, 
/* out0090_had-eta10-phi4*/	2, 66, 1, 67, 3, 
/* out0091_had-eta11-phi4*/	2, 66, 4, 123, 1, 
/* out0092_had-eta12-phi4*/	2, 66, 3, 123, 5, 
/* out0093_had-eta13-phi4*/	4, 60, 1, 89, 2, 121, 1, 123, 3, 
/* out0094_had-eta14-phi4*/	4, 60, 1, 89, 1, 116, 1, 121, 2, 
/* out0095_had-eta15-phi4*/	3, 88, 2, 120, 2, 121, 1, 
/* out0096_had-eta16-phi4*/	2, 88, 2, 120, 2, 
/* out0097_had-eta17-phi4*/	2, 88, 1, 120, 2, 
/* out0098_had-eta18-phi4*/	2, 88, 1, 120, 1, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	1, 143, 3, 
/* out0101_had-eta1-phi5*/	1, 143, 4, 
/* out0102_had-eta2-phi5*/	2, 142, 4, 143, 1, 
/* out0103_had-eta3-phi5*/	1, 142, 4, 
/* out0104_had-eta4-phi5*/	1, 141, 4, 
/* out0105_had-eta5-phi5*/	2, 74, 7, 141, 4, 
/* out0106_had-eta6-phi5*/	4, 72, 1, 74, 5, 77, 3, 140, 3, 
/* out0107_had-eta7-phi5*/	4, 71, 2, 72, 1, 77, 4, 140, 3, 
/* out0108_had-eta8-phi5*/	2, 71, 6, 140, 2, 
/* out0109_had-eta9-phi5*/	2, 71, 1, 75, 4, 
/* out0110_had-eta10-phi5*/	2, 66, 1, 75, 4, 
/* out0111_had-eta11-phi5*/	2, 66, 3, 123, 1, 
/* out0112_had-eta12-phi5*/	3, 60, 1, 66, 2, 123, 4, 
/* out0113_had-eta13-phi5*/	3, 60, 2, 116, 2, 123, 2, 
/* out0114_had-eta14-phi5*/	2, 60, 2, 116, 3, 
/* out0115_had-eta15-phi5*/	3, 60, 1, 88, 1, 116, 2, 
/* out0116_had-eta16-phi5*/	2, 88, 1, 120, 2, 
/* out0117_had-eta17-phi5*/	2, 88, 1, 120, 2, 
/* out0118_had-eta18-phi5*/	0, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	1, 147, 3, 
/* out0121_had-eta1-phi6*/	1, 147, 4, 
/* out0122_had-eta2-phi6*/	2, 146, 4, 147, 1, 
/* out0123_had-eta3-phi6*/	1, 146, 4, 
/* out0124_had-eta4-phi6*/	1, 145, 4, 
/* out0125_had-eta5-phi6*/	2, 79, 7, 145, 4, 
/* out0126_had-eta6-phi6*/	4, 77, 4, 78, 1, 79, 5, 144, 3, 
/* out0127_had-eta7-phi6*/	4, 76, 2, 77, 5, 78, 1, 144, 3, 
/* out0128_had-eta8-phi6*/	2, 76, 6, 144, 2, 
/* out0129_had-eta9-phi6*/	2, 75, 4, 76, 1, 
/* out0130_had-eta10-phi6*/	2, 61, 1, 75, 4, 
/* out0131_had-eta11-phi6*/	2, 61, 3, 118, 1, 
/* out0132_had-eta12-phi6*/	3, 60, 1, 61, 2, 118, 4, 
/* out0133_had-eta13-phi6*/	3, 60, 2, 116, 2, 118, 2, 
/* out0134_had-eta14-phi6*/	2, 60, 2, 116, 3, 
/* out0135_had-eta15-phi6*/	3, 53, 1, 60, 1, 116, 2, 
/* out0136_had-eta16-phi6*/	2, 53, 1, 115, 2, 
/* out0137_had-eta17-phi6*/	2, 53, 1, 115, 2, 
/* out0138_had-eta18-phi6*/	0, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	1, 147, 3, 
/* out0141_had-eta1-phi7*/	1, 147, 4, 
/* out0142_had-eta2-phi7*/	2, 146, 4, 147, 1, 
/* out0143_had-eta3-phi7*/	1, 146, 4, 
/* out0144_had-eta4-phi7*/	1, 145, 4, 
/* out0145_had-eta5-phi7*/	3, 79, 2, 80, 6, 145, 4, 
/* out0146_had-eta6-phi7*/	4, 78, 6, 79, 2, 80, 2, 144, 3, 
/* out0147_had-eta7-phi7*/	4, 63, 1, 76, 1, 78, 6, 144, 3, 
/* out0148_had-eta8-phi7*/	3, 63, 2, 76, 5, 144, 2, 
/* out0149_had-eta9-phi7*/	2, 62, 5, 76, 1, 
/* out0150_had-eta10-phi7*/	2, 61, 1, 62, 3, 
/* out0151_had-eta11-phi7*/	2, 61, 4, 118, 1, 
/* out0152_had-eta12-phi7*/	2, 61, 3, 118, 5, 
/* out0153_had-eta13-phi7*/	4, 54, 2, 60, 1, 117, 1, 118, 3, 
/* out0154_had-eta14-phi7*/	4, 54, 1, 60, 1, 116, 1, 117, 2, 
/* out0155_had-eta15-phi7*/	3, 53, 2, 115, 2, 117, 1, 
/* out0156_had-eta16-phi7*/	2, 53, 2, 115, 2, 
/* out0157_had-eta17-phi7*/	2, 53, 1, 115, 2, 
/* out0158_had-eta18-phi7*/	2, 53, 1, 115, 1, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	1, 151, 3, 
/* out0161_had-eta1-phi8*/	1, 151, 4, 
/* out0162_had-eta2-phi8*/	2, 150, 4, 151, 1, 
/* out0163_had-eta3-phi8*/	1, 150, 4, 
/* out0164_had-eta4-phi8*/	1, 149, 4, 
/* out0165_had-eta5-phi8*/	3, 65, 3, 80, 6, 149, 4, 
/* out0166_had-eta6-phi8*/	4, 64, 6, 78, 1, 80, 2, 148, 3, 
/* out0167_had-eta7-phi8*/	4, 63, 4, 64, 2, 78, 1, 148, 3, 
/* out0168_had-eta8-phi8*/	2, 63, 6, 148, 2, 
/* out0169_had-eta9-phi8*/	2, 56, 1, 62, 5, 
/* out0170_had-eta10-phi8*/	2, 55, 1, 62, 3, 
/* out0171_had-eta11-phi8*/	3, 55, 3, 61, 1, 119, 3, 
/* out0172_had-eta12-phi8*/	4, 54, 2, 55, 1, 61, 1, 119, 4, 
/* out0173_had-eta13-phi8*/	3, 54, 3, 117, 3, 119, 1, 
/* out0174_had-eta14-phi8*/	2, 54, 2, 117, 3, 
/* out0175_had-eta15-phi8*/	3, 53, 2, 115, 1, 117, 2, 
/* out0176_had-eta16-phi8*/	2, 53, 2, 115, 2, 
/* out0177_had-eta17-phi8*/	2, 53, 1, 115, 2, 
/* out0178_had-eta18-phi8*/	2, 46, 1, 111, 2, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	1, 151, 3, 
/* out0181_had-eta1-phi9*/	1, 151, 4, 
/* out0182_had-eta2-phi9*/	2, 150, 4, 151, 1, 
/* out0183_had-eta3-phi9*/	1, 150, 4, 
/* out0184_had-eta4-phi9*/	1, 149, 4, 
/* out0185_had-eta5-phi9*/	4, 58, 1, 59, 1, 65, 12, 149, 4, 
/* out0186_had-eta6-phi9*/	4, 58, 3, 64, 6, 65, 1, 148, 3, 
/* out0187_had-eta7-phi9*/	4, 57, 5, 63, 1, 64, 2, 148, 3, 
/* out0188_had-eta8-phi9*/	4, 56, 3, 57, 2, 63, 2, 148, 2, 
/* out0189_had-eta9-phi9*/	1, 56, 5, 
/* out0190_had-eta10-phi9*/	2, 55, 3, 56, 1, 
/* out0191_had-eta11-phi9*/	2, 55, 4, 119, 3, 
/* out0192_had-eta12-phi9*/	3, 54, 1, 55, 1, 119, 4, 
/* out0193_had-eta13-phi9*/	4, 54, 3, 113, 2, 117, 1, 119, 1, 
/* out0194_had-eta14-phi9*/	3, 54, 2, 113, 1, 117, 2, 
/* out0195_had-eta15-phi9*/	3, 47, 1, 112, 2, 117, 1, 
/* out0196_had-eta16-phi9*/	3, 47, 1, 53, 1, 112, 2, 
/* out0197_had-eta17-phi9*/	4, 46, 1, 53, 1, 111, 2, 112, 1, 
/* out0198_had-eta18-phi9*/	2, 46, 2, 111, 3, 
/* out0199_had-eta19-phi9*/	1, 111, 1, 
/* out0200_had-eta0-phi10*/	1, 155, 3, 
/* out0201_had-eta1-phi10*/	1, 155, 4, 
/* out0202_had-eta2-phi10*/	2, 154, 4, 155, 1, 
/* out0203_had-eta3-phi10*/	1, 154, 4, 
/* out0204_had-eta4-phi10*/	1, 153, 4, 
/* out0205_had-eta5-phi10*/	4, 52, 1, 58, 3, 59, 14, 153, 4, 
/* out0206_had-eta6-phi10*/	2, 58, 9, 152, 3, 
/* out0207_had-eta7-phi10*/	3, 51, 1, 57, 7, 152, 3, 
/* out0208_had-eta8-phi10*/	4, 50, 2, 56, 1, 57, 2, 152, 2, 
/* out0209_had-eta9-phi10*/	3, 49, 1, 50, 1, 56, 4, 
/* out0210_had-eta10-phi10*/	3, 49, 3, 55, 1, 56, 1, 
/* out0211_had-eta11-phi10*/	4, 48, 1, 49, 1, 55, 2, 114, 4, 
/* out0212_had-eta12-phi10*/	3, 48, 3, 113, 2, 114, 5, 
/* out0213_had-eta13-phi10*/	2, 48, 2, 113, 4, 
/* out0214_had-eta14-phi10*/	3, 47, 2, 112, 1, 113, 2, 
/* out0215_had-eta15-phi10*/	2, 47, 2, 112, 3, 
/* out0216_had-eta16-phi10*/	2, 47, 2, 112, 2, 
/* out0217_had-eta17-phi10*/	3, 46, 2, 111, 1, 112, 1, 
/* out0218_had-eta18-phi10*/	2, 46, 2, 111, 3, 
/* out0219_had-eta19-phi10*/	1, 111, 1, 
/* out0220_had-eta0-phi11*/	1, 155, 3, 
/* out0221_had-eta1-phi11*/	1, 155, 4, 
/* out0222_had-eta2-phi11*/	2, 154, 4, 155, 1, 
/* out0223_had-eta3-phi11*/	1, 154, 4, 
/* out0224_had-eta4-phi11*/	1, 153, 4, 
/* out0225_had-eta5-phi11*/	3, 52, 9, 59, 1, 153, 4, 
/* out0226_had-eta6-phi11*/	3, 51, 5, 52, 4, 152, 3, 
/* out0227_had-eta7-phi11*/	3, 50, 1, 51, 7, 152, 3, 
/* out0228_had-eta8-phi11*/	2, 50, 6, 152, 2, 
/* out0229_had-eta9-phi11*/	2, 49, 2, 50, 3, 
/* out0230_had-eta10-phi11*/	1, 49, 5, 
/* out0231_had-eta11-phi11*/	3, 48, 1, 49, 2, 114, 3, 
/* out0232_had-eta12-phi11*/	4, 48, 3, 110, 2, 113, 1, 114, 4, 
/* out0233_had-eta13-phi11*/	3, 48, 3, 110, 1, 113, 3, 
/* out0234_had-eta14-phi11*/	3, 47, 2, 109, 1, 113, 1, 
/* out0235_had-eta15-phi11*/	3, 47, 2, 109, 1, 112, 2, 
/* out0236_had-eta16-phi11*/	2, 47, 2, 112, 2, 
/* out0237_had-eta17-phi11*/	2, 46, 2, 108, 1, 
/* out0238_had-eta18-phi11*/	3, 46, 2, 108, 1, 111, 2, 
/* out0239_had-eta19-phi11*/	2, 46, 1, 111, 1, 
/* out0240_had-eta0-phi12*/	1, 159, 3, 
/* out0241_had-eta1-phi12*/	1, 159, 4, 
/* out0242_had-eta2-phi12*/	2, 158, 4, 159, 1, 
/* out0243_had-eta3-phi12*/	1, 158, 4, 
/* out0244_had-eta4-phi12*/	1, 157, 4, 
/* out0245_had-eta5-phi12*/	4, 44, 2, 45, 11, 52, 2, 157, 4, 
/* out0246_had-eta6-phi12*/	3, 44, 8, 51, 1, 156, 3, 
/* out0247_had-eta7-phi12*/	3, 43, 5, 51, 2, 156, 3, 
/* out0248_had-eta8-phi12*/	4, 42, 1, 43, 3, 50, 2, 156, 2, 
/* out0249_had-eta9-phi12*/	2, 42, 5, 50, 1, 
/* out0250_had-eta10-phi12*/	3, 41, 1, 42, 1, 49, 2, 
/* out0251_had-eta11-phi12*/	2, 41, 3, 110, 2, 
/* out0252_had-eta12-phi12*/	3, 41, 1, 48, 2, 110, 4, 
/* out0253_had-eta13-phi12*/	4, 40, 2, 48, 1, 109, 1, 110, 3, 
/* out0254_had-eta14-phi12*/	2, 40, 2, 109, 3, 
/* out0255_had-eta15-phi12*/	2, 47, 1, 109, 3, 
/* out0256_had-eta16-phi12*/	4, 39, 1, 47, 1, 108, 2, 109, 1, 
/* out0257_had-eta17-phi12*/	2, 39, 1, 108, 2, 
/* out0258_had-eta18-phi12*/	2, 46, 2, 108, 2, 
/* out0259_had-eta19-phi12*/	2, 46, 1, 108, 1, 
/* out0260_had-eta0-phi13*/	1, 159, 3, 
/* out0261_had-eta1-phi13*/	1, 159, 4, 
/* out0262_had-eta2-phi13*/	2, 158, 4, 159, 1, 
/* out0263_had-eta3-phi13*/	1, 158, 4, 
/* out0264_had-eta4-phi13*/	1, 157, 4, 
/* out0265_had-eta5-phi13*/	4, 38, 8, 44, 1, 45, 5, 157, 4, 
/* out0266_had-eta6-phi13*/	4, 37, 3, 38, 1, 44, 5, 156, 3, 
/* out0267_had-eta7-phi13*/	3, 37, 3, 43, 5, 156, 3, 
/* out0268_had-eta8-phi13*/	4, 36, 2, 42, 2, 43, 3, 156, 2, 
/* out0269_had-eta9-phi13*/	1, 42, 5, 
/* out0270_had-eta10-phi13*/	2, 41, 2, 42, 2, 
/* out0271_had-eta11-phi13*/	2, 41, 4, 107, 3, 
/* out0272_had-eta12-phi13*/	4, 40, 1, 41, 2, 107, 2, 110, 3, 
/* out0273_had-eta13-phi13*/	4, 40, 3, 105, 2, 109, 1, 110, 1, 
/* out0274_had-eta14-phi13*/	2, 40, 2, 109, 3, 
/* out0275_had-eta15-phi13*/	3, 39, 1, 40, 1, 109, 2, 
/* out0276_had-eta16-phi13*/	2, 39, 2, 108, 2, 
/* out0277_had-eta17-phi13*/	2, 39, 1, 108, 2, 
/* out0278_had-eta18-phi13*/	2, 39, 1, 108, 1, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	1, 163, 3, 
/* out0281_had-eta1-phi14*/	1, 163, 4, 
/* out0282_had-eta2-phi14*/	2, 162, 4, 163, 1, 
/* out0283_had-eta3-phi14*/	1, 162, 4, 
/* out0284_had-eta4-phi14*/	1, 161, 4, 
/* out0285_had-eta5-phi14*/	3, 32, 3, 38, 6, 161, 4, 
/* out0286_had-eta6-phi14*/	4, 32, 2, 37, 6, 38, 1, 160, 3, 
/* out0287_had-eta7-phi14*/	4, 31, 1, 36, 3, 37, 4, 160, 3, 
/* out0288_had-eta8-phi14*/	2, 36, 7, 160, 2, 
/* out0289_had-eta9-phi14*/	2, 35, 4, 36, 2, 
/* out0290_had-eta10-phi14*/	1, 35, 4, 
/* out0291_had-eta11-phi14*/	4, 34, 1, 35, 1, 41, 2, 107, 6, 
/* out0292_had-eta12-phi14*/	4, 34, 2, 41, 1, 105, 3, 107, 4, 
/* out0293_had-eta13-phi14*/	2, 40, 2, 105, 4, 
/* out0294_had-eta14-phi14*/	3, 40, 2, 103, 1, 105, 2, 
/* out0295_had-eta15-phi14*/	3, 39, 1, 40, 1, 103, 3, 
/* out0296_had-eta16-phi14*/	2, 39, 2, 103, 2, 
/* out0297_had-eta17-phi14*/	2, 39, 1, 108, 1, 
/* out0298_had-eta18-phi14*/	3, 39, 1, 102, 1, 108, 1, 
/* out0299_had-eta19-phi14*/	1, 102, 1, 
/* out0300_had-eta0-phi15*/	1, 163, 3, 
/* out0301_had-eta1-phi15*/	1, 163, 4, 
/* out0302_had-eta2-phi15*/	2, 162, 4, 163, 1, 
/* out0303_had-eta3-phi15*/	1, 162, 4, 
/* out0304_had-eta4-phi15*/	1, 161, 4, 
/* out0305_had-eta5-phi15*/	3, 28, 7, 32, 6, 161, 4, 
/* out0306_had-eta6-phi15*/	4, 26, 1, 31, 3, 32, 5, 160, 3, 
/* out0307_had-eta7-phi15*/	2, 31, 8, 160, 3, 
/* out0308_had-eta8-phi15*/	3, 30, 4, 36, 2, 160, 2, 
/* out0309_had-eta9-phi15*/	2, 30, 2, 35, 3, 
/* out0310_had-eta10-phi15*/	1, 35, 4, 
/* out0311_had-eta11-phi15*/	3, 34, 4, 106, 4, 107, 1, 
/* out0312_had-eta12-phi15*/	3, 34, 3, 105, 1, 106, 4, 
/* out0313_had-eta13-phi15*/	4, 33, 1, 34, 1, 104, 1, 105, 3, 
/* out0314_had-eta14-phi15*/	4, 33, 2, 103, 2, 104, 1, 105, 1, 
/* out0315_had-eta15-phi15*/	2, 33, 1, 103, 3, 
/* out0316_had-eta16-phi15*/	2, 39, 2, 103, 2, 
/* out0317_had-eta17-phi15*/	2, 39, 1, 102, 2, 
/* out0318_had-eta18-phi15*/	2, 39, 1, 102, 2, 
/* out0319_had-eta19-phi15*/	1, 102, 1, 
/* out0320_had-eta0-phi16*/	1, 167, 3, 
/* out0321_had-eta1-phi16*/	1, 167, 4, 
/* out0322_had-eta2-phi16*/	2, 166, 4, 167, 1, 
/* out0323_had-eta3-phi16*/	1, 166, 4, 
/* out0324_had-eta4-phi16*/	1, 165, 4, 
/* out0325_had-eta5-phi16*/	4, 26, 4, 27, 3, 28, 9, 165, 4, 
/* out0326_had-eta6-phi16*/	3, 26, 8, 31, 1, 164, 3, 
/* out0327_had-eta7-phi16*/	3, 25, 5, 31, 3, 164, 3, 
/* out0328_had-eta8-phi16*/	3, 25, 1, 30, 6, 164, 2, 
/* out0329_had-eta9-phi16*/	2, 29, 2, 30, 4, 
/* out0330_had-eta10-phi16*/	1, 29, 4, 
/* out0331_had-eta11-phi16*/	3, 29, 2, 34, 2, 106, 3, 
/* out0332_had-eta12-phi16*/	4, 14, 1, 34, 2, 104, 1, 106, 5, 
/* out0333_had-eta13-phi16*/	3, 33, 2, 34, 1, 104, 4, 
/* out0334_had-eta14-phi16*/	2, 33, 2, 104, 3, 
/* out0335_had-eta15-phi16*/	3, 33, 2, 98, 1, 103, 2, 
/* out0336_had-eta16-phi16*/	4, 0, 1, 33, 1, 98, 1, 103, 1, 
/* out0337_had-eta17-phi16*/	2, 0, 1, 102, 2, 
/* out0338_had-eta18-phi16*/	2, 0, 1, 102, 2, 
/* out0339_had-eta19-phi16*/	1, 102, 1, 
/* out0340_had-eta0-phi17*/	1, 167, 3, 
/* out0341_had-eta1-phi17*/	1, 167, 4, 
/* out0342_had-eta2-phi17*/	2, 166, 4, 167, 1, 
/* out0343_had-eta3-phi17*/	1, 166, 4, 
/* out0344_had-eta4-phi17*/	1, 165, 4, 
/* out0345_had-eta5-phi17*/	4, 23, 2, 26, 1, 27, 13, 165, 4, 
/* out0346_had-eta6-phi17*/	4, 23, 6, 25, 1, 26, 2, 164, 3, 
/* out0347_had-eta7-phi17*/	2, 25, 8, 164, 3, 
/* out0348_had-eta8-phi17*/	3, 19, 4, 25, 1, 164, 2, 
/* out0349_had-eta9-phi17*/	2, 19, 3, 29, 2, 
/* out0350_had-eta10-phi17*/	1, 29, 4, 
/* out0351_had-eta11-phi17*/	3, 14, 2, 29, 2, 101, 3, 
/* out0352_had-eta12-phi17*/	2, 14, 3, 101, 5, 
/* out0353_had-eta13-phi17*/	3, 14, 2, 33, 1, 104, 3, 
/* out0354_had-eta14-phi17*/	2, 33, 2, 104, 3, 
/* out0355_had-eta15-phi17*/	2, 33, 2, 98, 3, 
/* out0356_had-eta16-phi17*/	2, 0, 2, 98, 2, 
/* out0357_had-eta17-phi17*/	3, 0, 2, 98, 1, 102, 1, 
/* out0358_had-eta18-phi17*/	2, 0, 1, 102, 2, 
/* out0359_had-eta19-phi17*/	1, 102, 1, 
/* out0360_had-eta0-phi18*/	1, 171, 3, 
/* out0361_had-eta1-phi18*/	1, 171, 4, 
/* out0362_had-eta2-phi18*/	2, 170, 4, 171, 1, 
/* out0363_had-eta3-phi18*/	1, 170, 4, 
/* out0364_had-eta4-phi18*/	1, 169, 4, 
/* out0365_had-eta5-phi18*/	4, 21, 1, 23, 2, 24, 13, 169, 4, 
/* out0366_had-eta6-phi18*/	4, 20, 1, 21, 2, 23, 6, 168, 3, 
/* out0367_had-eta7-phi18*/	2, 20, 8, 168, 3, 
/* out0368_had-eta8-phi18*/	3, 19, 5, 20, 1, 168, 2, 
/* out0369_had-eta9-phi18*/	2, 15, 2, 19, 4, 
/* out0370_had-eta10-phi18*/	1, 15, 4, 
/* out0371_had-eta11-phi18*/	3, 14, 2, 15, 2, 101, 3, 
/* out0372_had-eta12-phi18*/	2, 14, 3, 101, 5, 
/* out0373_had-eta13-phi18*/	3, 1, 1, 14, 2, 99, 3, 
/* out0374_had-eta14-phi18*/	2, 1, 2, 99, 3, 
/* out0375_had-eta15-phi18*/	2, 1, 2, 98, 3, 
/* out0376_had-eta16-phi18*/	2, 0, 2, 98, 2, 
/* out0377_had-eta17-phi18*/	3, 0, 2, 98, 1, 128, 1, 
/* out0378_had-eta18-phi18*/	2, 0, 1, 128, 2, 
/* out0379_had-eta19-phi18*/	1, 128, 1, 
/* out0380_had-eta0-phi19*/	1, 171, 3, 
/* out0381_had-eta1-phi19*/	1, 171, 4, 
/* out0382_had-eta2-phi19*/	2, 170, 4, 171, 1, 
/* out0383_had-eta3-phi19*/	1, 170, 4, 
/* out0384_had-eta4-phi19*/	1, 169, 4, 
/* out0385_had-eta5-phi19*/	4, 21, 4, 22, 9, 24, 3, 169, 4, 
/* out0386_had-eta6-phi19*/	3, 17, 1, 21, 8, 168, 3, 
/* out0387_had-eta7-phi19*/	3, 17, 3, 20, 5, 168, 3, 
/* out0388_had-eta8-phi19*/	3, 16, 6, 20, 1, 168, 2, 
/* out0389_had-eta9-phi19*/	2, 15, 2, 16, 4, 
/* out0390_had-eta10-phi19*/	1, 15, 4, 
/* out0391_had-eta11-phi19*/	3, 2, 2, 15, 2, 100, 3, 
/* out0392_had-eta12-phi19*/	4, 2, 2, 14, 1, 99, 1, 100, 5, 
/* out0393_had-eta13-phi19*/	3, 1, 2, 2, 1, 99, 4, 
/* out0394_had-eta14-phi19*/	2, 1, 2, 99, 3, 
/* out0395_had-eta15-phi19*/	3, 1, 2, 98, 1, 129, 2, 
/* out0396_had-eta16-phi19*/	4, 0, 1, 1, 1, 98, 1, 129, 1, 
/* out0397_had-eta17-phi19*/	2, 0, 1, 128, 2, 
/* out0398_had-eta18-phi19*/	2, 0, 1, 128, 2, 
/* out0399_had-eta19-phi19*/	1, 128, 1, 
/* out0400_had-eta0-phi20*/	1, 175, 3, 
/* out0401_had-eta1-phi20*/	1, 175, 4, 
/* out0402_had-eta2-phi20*/	2, 174, 4, 175, 1, 
/* out0403_had-eta3-phi20*/	1, 174, 4, 
/* out0404_had-eta4-phi20*/	1, 173, 4, 
/* out0405_had-eta5-phi20*/	3, 18, 6, 22, 7, 173, 4, 
/* out0406_had-eta6-phi20*/	4, 17, 3, 18, 5, 21, 1, 172, 3, 
/* out0407_had-eta7-phi20*/	2, 17, 8, 172, 3, 
/* out0408_had-eta8-phi20*/	3, 4, 2, 16, 4, 172, 2, 
/* out0409_had-eta9-phi20*/	2, 3, 3, 16, 2, 
/* out0410_had-eta10-phi20*/	1, 3, 4, 
/* out0411_had-eta11-phi20*/	3, 2, 4, 100, 4, 131, 1, 
/* out0412_had-eta12-phi20*/	3, 2, 3, 100, 4, 130, 1, 
/* out0413_had-eta13-phi20*/	4, 1, 1, 2, 1, 99, 1, 130, 3, 
/* out0414_had-eta14-phi20*/	4, 1, 2, 99, 1, 129, 2, 130, 1, 
/* out0415_had-eta15-phi20*/	2, 1, 1, 129, 3, 
/* out0416_had-eta16-phi20*/	2, 7, 2, 129, 2, 
/* out0417_had-eta17-phi20*/	2, 7, 1, 128, 2, 
/* out0418_had-eta18-phi20*/	2, 7, 1, 128, 2, 
/* out0419_had-eta19-phi20*/	1, 128, 1, 
/* out0420_had-eta0-phi21*/	1, 175, 3, 
/* out0421_had-eta1-phi21*/	1, 175, 4, 
/* out0422_had-eta2-phi21*/	2, 174, 4, 175, 1, 
/* out0423_had-eta3-phi21*/	1, 174, 4, 
/* out0424_had-eta4-phi21*/	1, 173, 4, 
/* out0425_had-eta5-phi21*/	3, 6, 6, 18, 3, 173, 4, 
/* out0426_had-eta6-phi21*/	4, 5, 6, 6, 1, 18, 2, 172, 3, 
/* out0427_had-eta7-phi21*/	4, 4, 3, 5, 4, 17, 1, 172, 3, 
/* out0428_had-eta8-phi21*/	2, 4, 7, 172, 2, 
/* out0429_had-eta9-phi21*/	2, 3, 4, 4, 2, 
/* out0430_had-eta10-phi21*/	1, 3, 4, 
/* out0431_had-eta11-phi21*/	4, 2, 1, 3, 1, 9, 2, 131, 6, 
/* out0432_had-eta12-phi21*/	4, 2, 2, 9, 1, 130, 3, 131, 4, 
/* out0433_had-eta13-phi21*/	2, 8, 2, 130, 4, 
/* out0434_had-eta14-phi21*/	3, 8, 2, 129, 1, 130, 2, 
/* out0435_had-eta15-phi21*/	3, 7, 1, 8, 1, 129, 3, 
/* out0436_had-eta16-phi21*/	2, 7, 2, 129, 2, 
/* out0437_had-eta17-phi21*/	2, 7, 1, 95, 1, 
/* out0438_had-eta18-phi21*/	3, 7, 1, 95, 1, 128, 1, 
/* out0439_had-eta19-phi21*/	1, 128, 1, 
/* out0440_had-eta0-phi22*/	1, 179, 3, 
/* out0441_had-eta1-phi22*/	1, 179, 4, 
/* out0442_had-eta2-phi22*/	2, 178, 4, 179, 1, 
/* out0443_had-eta3-phi22*/	1, 178, 4, 
/* out0444_had-eta4-phi22*/	1, 177, 4, 
/* out0445_had-eta5-phi22*/	4, 6, 8, 12, 1, 13, 5, 177, 4, 
/* out0446_had-eta6-phi22*/	4, 5, 3, 6, 1, 12, 5, 176, 3, 
/* out0447_had-eta7-phi22*/	3, 5, 3, 11, 5, 176, 3, 
/* out0448_had-eta8-phi22*/	4, 4, 2, 10, 2, 11, 3, 176, 2, 
/* out0449_had-eta9-phi22*/	1, 10, 5, 
/* out0450_had-eta10-phi22*/	2, 9, 2, 10, 2, 
/* out0451_had-eta11-phi22*/	3, 9, 4, 97, 1, 131, 3, 
/* out0452_had-eta12-phi22*/	4, 8, 1, 9, 2, 97, 3, 131, 2, 
/* out0453_had-eta13-phi22*/	4, 8, 3, 96, 1, 97, 2, 130, 2, 
/* out0454_had-eta14-phi22*/	2, 8, 2, 96, 3, 
/* out0455_had-eta15-phi22*/	3, 7, 1, 8, 1, 96, 3, 
/* out0456_had-eta16-phi22*/	2, 7, 2, 95, 2, 
/* out0457_had-eta17-phi22*/	2, 7, 1, 95, 2, 
/* out0458_had-eta18-phi22*/	2, 7, 1, 95, 2, 
/* out0459_had-eta19-phi22*/	1, 95, 1, 
/* out0460_had-eta0-phi23*/	1, 179, 3, 
/* out0461_had-eta1-phi23*/	1, 179, 4, 
/* out0462_had-eta2-phi23*/	2, 178, 4, 179, 1, 
/* out0463_had-eta3-phi23*/	1, 178, 4, 
/* out0464_had-eta4-phi23*/	1, 177, 4, 
/* out0465_had-eta5-phi23*/	3, 12, 2, 13, 11, 177, 4, 
/* out0466_had-eta6-phi23*/	2, 12, 8, 176, 3, 
/* out0467_had-eta7-phi23*/	2, 11, 5, 176, 3, 
/* out0468_had-eta8-phi23*/	3, 10, 1, 11, 3, 176, 2, 
/* out0469_had-eta9-phi23*/	1, 10, 5, 
/* out0470_had-eta10-phi23*/	2, 9, 1, 10, 1, 
/* out0471_had-eta11-phi23*/	2, 9, 3, 97, 2, 
/* out0472_had-eta12-phi23*/	2, 9, 1, 97, 5, 
/* out0473_had-eta13-phi23*/	3, 8, 2, 96, 1, 97, 3, 
/* out0474_had-eta14-phi23*/	2, 8, 2, 96, 4, 
/* out0475_had-eta15-phi23*/	1, 96, 3, 
/* out0476_had-eta16-phi23*/	3, 7, 1, 95, 2, 96, 1, 
/* out0477_had-eta17-phi23*/	2, 7, 1, 95, 2, 
/* out0478_had-eta18-phi23*/	1, 95, 2, 
/* out0479_had-eta19-phi23*/	1, 95, 1, 
};