parameter integer matrixH [0:7775] = {
/* num inputs = 133(in0-in132) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2431 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	1,110,0,14,
/* out0002_em-eta2-phi0*/	2,110,0,2,110,1,16,
/* out0003_em-eta3-phi0*/	2,109,0,16,109,1,2,
/* out0004_em-eta4-phi0*/	2,87,2,2,109,1,14,
/* out0005_em-eta5-phi0*/	4,86,0,3,86,1,6,87,1,8,87,2,13,
/* out0006_em-eta6-phi0*/	7,58,2,1,63,0,1,63,1,6,85,1,1,86,0,13,86,1,2,86,2,7,
/* out0007_em-eta7-phi0*/	6,63,0,8,63,1,8,63,2,9,85,0,13,85,1,4,85,2,1,
/* out0008_em-eta8-phi0*/	8,62,0,4,62,1,12,63,0,7,63,2,4,84,0,3,84,1,3,85,0,3,85,2,3,
/* out0009_em-eta9-phi0*/	6,61,0,7,61,1,1,62,0,12,62,2,11,84,0,12,84,2,1,
/* out0010_em-eta10-phi0*/	7,61,0,5,61,1,9,61,2,1,83,0,3,83,1,1,84,0,1,84,2,1,
/* out0011_em-eta11-phi0*/	7,60,0,6,60,1,1,61,0,4,61,2,8,104,0,2,104,1,6,83,0,9,
/* out0012_em-eta12-phi0*/	8,60,0,4,60,1,7,104,0,7,104,1,3,104,2,4,82,0,1,82,1,1,83,0,2,
/* out0013_em-eta13-phi0*/	7,60,0,5,60,2,3,103,0,1,103,1,4,104,0,7,104,2,5,82,0,6,
/* out0014_em-eta14-phi0*/	8,59,0,1,59,1,3,60,0,1,60,2,3,103,0,6,103,1,3,103,2,1,82,0,4,
/* out0015_em-eta15-phi0*/	5,59,0,4,59,1,2,103,0,3,103,2,5,81,0,1,
/* out0016_em-eta16-phi0*/	6,59,0,10,59,2,2,102,0,2,102,1,4,103,0,6,81,0,3,
/* out0017_em-eta17-phi0*/	5,59,0,1,59,2,2,102,0,5,102,1,1,81,0,3,
/* out0018_em-eta18-phi0*/	2,102,0,8,102,2,2,
/* out0019_em-eta19-phi0*/	2,102,0,1,102,2,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	1,110,3,14,
/* out0022_em-eta2-phi1*/	2,110,2,16,110,3,2,
/* out0023_em-eta3-phi1*/	2,109,2,2,109,3,16,
/* out0024_em-eta4-phi1*/	4,80,1,3,87,1,1,87,2,1,109,2,14,
/* out0025_em-eta5-phi1*/	5,80,0,16,80,1,4,80,2,3,86,1,5,87,1,7,
/* out0026_em-eta6-phi1*/	8,58,1,2,58,2,10,79,0,10,79,1,2,80,2,1,85,1,1,86,1,3,86,2,9,
/* out0027_em-eta7-phi1*/	10,57,0,5,57,1,7,58,1,7,58,2,4,63,1,2,63,2,3,78,0,2,79,0,4,85,1,10,85,2,7,
/* out0028_em-eta8-phi1*/	7,56,1,1,57,0,11,57,2,5,62,1,4,78,0,6,84,1,8,85,2,5,
/* out0029_em-eta9-phi1*/	5,56,0,10,56,1,2,62,2,5,84,1,5,84,2,10,
/* out0030_em-eta10-phi1*/	8,55,0,1,56,0,5,56,2,1,61,1,6,61,2,2,77,0,1,83,1,9,84,2,3,
/* out0031_em-eta11-phi1*/	7,55,0,6,61,2,5,100,2,9,104,1,3,83,0,2,83,1,3,83,2,6,
/* out0032_em-eta12-phi1*/	8,55,0,2,60,1,8,98,0,3,100,2,1,104,1,4,104,2,5,82,1,4,83,2,5,
/* out0033_em-eta13-phi1*/	7,60,2,8,98,0,6,103,1,3,104,2,2,82,0,3,82,1,4,82,2,1,
/* out0034_em-eta14-phi1*/	7,54,0,1,59,1,4,60,2,2,103,1,6,103,2,3,82,0,2,82,2,4,
/* out0035_em-eta15-phi1*/	7,59,1,5,59,2,1,97,0,1,103,2,6,81,0,1,81,1,3,82,2,2,
/* out0036_em-eta16-phi1*/	5,59,2,5,97,0,1,102,1,6,81,0,3,81,1,1,
/* out0037_em-eta17-phi1*/	4,59,2,2,102,1,3,102,2,3,81,0,3,
/* out0038_em-eta18-phi1*/	3,102,2,5,81,0,2,81,2,1,
/* out0039_em-eta19-phi1*/	1,102,2,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	1,112,0,14,
/* out0042_em-eta2-phi2*/	2,112,0,2,112,1,16,
/* out0043_em-eta3-phi2*/	2,111,0,16,111,1,2,
/* out0044_em-eta4-phi2*/	2,80,1,2,111,1,14,
/* out0045_em-eta5-phi2*/	4,74,0,8,74,1,2,80,1,7,80,2,11,
/* out0046_em-eta6-phi2*/	9,51,0,7,51,2,4,58,1,5,58,2,1,74,0,4,79,0,2,79,1,14,79,2,7,80,2,1,
/* out0047_em-eta7-phi2*/	10,49,1,1,51,0,1,51,1,3,51,2,12,57,1,9,58,1,2,73,0,2,78,0,1,78,1,11,79,2,9,
/* out0048_em-eta8-phi2*/	6,49,0,8,56,1,2,57,2,11,78,0,7,78,1,2,78,2,9,
/* out0049_em-eta9-phi2*/	8,49,0,1,56,0,1,56,1,11,56,2,5,77,0,6,77,1,7,78,2,1,84,2,1,
/* out0050_em-eta10-phi2*/	5,55,1,5,56,2,9,77,0,9,77,2,3,83,1,2,
/* out0051_em-eta11-phi2*/	9,55,0,4,55,1,6,55,2,2,100,1,10,100,2,6,76,0,4,76,1,1,83,1,1,83,2,4,
/* out0052_em-eta12-phi2*/	9,54,1,1,55,0,3,55,2,5,98,0,1,98,1,9,100,1,4,76,0,6,82,1,2,83,2,1,
/* out0053_em-eta13-phi2*/	7,54,0,5,54,1,3,98,0,5,98,1,1,98,2,5,82,1,5,82,2,2,
/* out0054_em-eta14-phi2*/	8,54,0,7,97,0,1,97,1,3,98,0,1,98,2,3,103,2,1,75,0,1,82,2,6,
/* out0055_em-eta15-phi2*/	8,53,1,1,54,0,2,59,1,2,59,2,1,97,0,7,97,1,1,81,1,4,82,2,1,
/* out0056_em-eta16-phi2*/	5,53,1,2,59,2,2,97,0,5,102,1,1,81,1,4,
/* out0057_em-eta17-phi2*/	7,53,0,1,53,1,1,59,2,1,96,1,1,102,1,1,102,2,2,81,2,4,
/* out0058_em-eta18-phi2*/	3,96,1,3,102,2,2,81,2,3,
/* out0059_em-eta19-phi2*/	1,96,0,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	1,112,3,14,
/* out0062_em-eta2-phi3*/	2,112,2,16,112,3,2,
/* out0063_em-eta3-phi3*/	2,111,2,2,111,3,16,
/* out0064_em-eta4-phi3*/	3,69,0,3,69,2,7,111,2,14,
/* out0065_em-eta5-phi3*/	7,68,0,1,69,0,1,69,1,8,69,2,9,74,0,2,74,1,14,74,2,7,
/* out0066_em-eta6-phi3*/	8,51,0,7,51,1,1,52,2,1,68,0,2,73,0,3,73,1,12,74,0,2,74,2,9,
/* out0067_em-eta7-phi3*/	9,49,1,5,51,0,1,51,1,12,52,1,6,72,1,1,73,0,11,73,1,1,73,2,8,78,1,2,
/* out0068_em-eta8-phi3*/	7,49,0,5,49,1,9,49,2,6,72,0,10,72,1,3,78,1,1,78,2,6,
/* out0069_em-eta9-phi3*/	8,48,0,3,48,1,6,49,0,2,49,2,5,56,2,1,72,0,4,77,1,9,77,2,3,
/* out0070_em-eta10-phi3*/	5,48,0,12,55,1,1,71,0,1,76,1,1,77,2,10,
/* out0071_em-eta11-phi3*/	10,47,0,2,48,0,1,48,2,1,55,1,4,55,2,5,100,1,2,101,0,8,101,2,9,76,0,1,76,1,10,
/* out0072_em-eta12-phi3*/	8,47,0,3,54,1,3,55,2,4,98,1,5,101,1,2,101,2,7,76,0,4,76,2,5,
/* out0073_em-eta13-phi3*/	9,54,1,7,54,2,1,98,1,1,98,2,7,99,1,3,75,0,1,75,1,3,76,0,1,76,2,2,
/* out0074_em-eta14-phi3*/	6,54,0,1,54,2,6,97,1,6,98,2,1,99,1,2,75,0,6,
/* out0075_em-eta15-phi3*/	7,53,1,3,54,2,3,97,0,1,97,1,4,97,2,3,75,0,4,81,1,1,
/* out0076_em-eta16-phi3*/	4,53,1,4,97,2,6,81,1,3,81,2,2,
/* out0077_em-eta17-phi3*/	4,53,0,5,53,1,1,96,1,5,81,2,4,
/* out0078_em-eta18-phi3*/	3,96,0,2,96,1,3,81,2,2,
/* out0079_em-eta19-phi3*/	1,96,0,3,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	1,114,0,14,
/* out0082_em-eta2-phi4*/	2,114,0,2,114,1,16,
/* out0083_em-eta3-phi4*/	2,113,0,16,113,1,2,
/* out0084_em-eta4-phi4*/	2,69,0,3,113,1,14,
/* out0085_em-eta5-phi4*/	7,68,0,3,68,1,14,68,2,1,69,0,9,69,1,8,70,0,5,70,1,6,
/* out0086_em-eta6-phi4*/	6,52,2,8,67,1,3,68,0,10,68,2,9,73,1,3,73,2,1,
/* out0087_em-eta7-phi4*/	7,52,0,10,52,1,9,52,2,6,67,0,12,67,1,1,72,1,3,73,2,7,
/* out0088_em-eta8-phi4*/	9,49,1,1,49,2,4,50,1,8,50,2,5,52,0,1,52,1,1,72,0,1,72,1,9,72,2,8,
/* out0089_em-eta9-phi4*/	8,48,1,9,48,2,1,49,2,1,50,1,7,71,0,1,71,1,7,72,0,1,72,2,7,
/* out0090_em-eta10-phi4*/	5,48,1,1,48,2,13,71,0,11,71,1,1,71,2,1,
/* out0091_em-eta11-phi4*/	10,47,0,2,47,1,9,48,2,1,101,0,8,101,1,6,56,1,1,71,0,3,71,2,1,76,1,4,76,2,2,
/* out0092_em-eta12-phi4*/	6,47,0,8,47,2,2,99,2,5,101,1,8,56,1,2,76,2,6,
/* out0093_em-eta13-phi4*/	10,42,1,1,47,0,1,47,2,1,54,1,2,54,2,2,99,0,1,99,1,5,99,2,5,75,1,7,76,2,1,
/* out0094_em-eta14-phi4*/	8,42,1,3,54,2,4,97,1,1,99,0,2,99,1,6,75,0,2,75,1,2,75,2,2,
/* out0095_em-eta15-phi4*/	8,42,1,1,53,1,2,53,2,3,92,1,2,97,1,1,97,2,4,75,0,2,75,2,4,
/* out0096_em-eta16-phi4*/	8,53,1,2,53,2,3,92,1,2,96,1,1,96,2,1,97,2,3,75,2,1,88,1,2,
/* out0097_em-eta17-phi4*/	4,53,0,7,96,1,2,96,2,3,88,1,3,
/* out0098_em-eta18-phi4*/	5,96,0,3,96,1,1,96,2,2,88,0,2,88,1,1,
/* out0099_em-eta19-phi4*/	1,96,0,4,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	1,114,3,14,
/* out0102_em-eta2-phi5*/	2,114,2,16,114,3,2,
/* out0103_em-eta3-phi5*/	2,113,2,2,113,3,16,
/* out0104_em-eta4-phi5*/	1,113,2,14,
/* out0105_em-eta5-phi5*/	7,63,0,2,63,1,7,68,1,2,68,2,2,70,0,11,70,1,10,70,2,16,
/* out0106_em-eta6-phi5*/	4,66,1,3,63,0,14,67,1,8,68,2,4,
/* out0107_em-eta7-phi5*/	8,50,2,1,52,0,5,52,2,1,66,0,14,66,1,5,67,0,3,67,1,4,67,2,15,
/* out0108_em-eta8-phi5*/	8,50,0,7,50,2,10,66,0,2,61,1,8,61,2,7,67,0,1,67,2,1,72,2,1,
/* out0109_em-eta9-phi5*/	6,50,0,9,50,1,1,64,1,1,64,2,6,61,1,8,71,1,6,
/* out0110_em-eta10-phi5*/	4,64,1,12,64,2,2,71,1,2,71,2,11,
/* out0111_em-eta11-phi5*/	8,47,1,7,47,2,2,64,1,3,94,0,9,94,2,5,56,1,1,56,2,7,71,2,3,
/* out0112_em-eta12-phi5*/	6,47,2,10,94,1,1,94,2,11,99,2,2,56,1,8,56,2,1,
/* out0113_em-eta13-phi5*/	7,42,1,1,42,2,6,47,2,1,99,0,7,99,2,4,56,1,4,75,1,3,
/* out0114_em-eta14-phi5*/	6,42,1,6,42,2,1,92,2,2,99,0,6,75,1,1,75,2,5,
/* out0115_em-eta15-phi5*/	6,42,1,4,53,2,1,92,1,3,92,2,5,75,2,4,88,1,1,
/* out0116_em-eta16-phi5*/	3,53,2,6,92,1,7,88,1,4,
/* out0117_em-eta17-phi5*/	6,53,0,2,53,2,3,92,1,2,96,2,4,88,0,1,88,1,3,
/* out0118_em-eta18-phi5*/	3,53,0,1,96,2,5,88,0,4,
/* out0119_em-eta19-phi5*/	2,96,0,3,96,2,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	1,116,0,14,
/* out0122_em-eta2-phi6*/	2,116,0,2,116,1,16,
/* out0123_em-eta3-phi6*/	2,115,0,16,115,1,2,
/* out0124_em-eta4-phi6*/	1,115,1,14,
/* out0125_em-eta5-phi6*/	7,63,1,8,63,2,2,64,1,2,64,2,2,65,0,11,65,1,14,65,2,16,
/* out0126_em-eta6-phi6*/	5,66,1,3,62,2,8,63,1,1,63,2,14,64,1,4,
/* out0127_em-eta7-phi6*/	9,65,2,1,66,1,5,66,2,14,67,1,5,67,2,1,61,2,1,62,0,3,62,1,15,62,2,4,
/* out0128_em-eta8-phi6*/	8,65,1,7,65,2,10,66,2,2,58,1,1,61,0,8,61,2,8,62,0,1,62,1,1,
/* out0129_em-eta9-phi6*/	6,64,0,1,64,2,6,65,0,1,65,1,9,57,2,6,61,0,8,
/* out0130_em-eta10-phi6*/	4,64,0,12,64,2,2,57,1,11,57,2,2,
/* out0131_em-eta11-phi6*/	8,43,1,2,43,2,7,64,0,3,94,0,7,94,1,5,56,0,1,56,2,7,57,1,3,
/* out0132_em-eta12-phi6*/	5,43,1,10,93,2,2,94,1,10,56,0,8,56,2,1,
/* out0133_em-eta13-phi6*/	6,42,2,7,43,1,1,93,1,7,93,2,4,56,0,4,89,2,3,
/* out0134_em-eta14-phi6*/	6,42,0,6,42,2,1,92,2,3,93,1,6,89,1,5,89,2,1,
/* out0135_em-eta15-phi6*/	6,36,1,1,42,0,5,92,0,3,92,2,5,88,2,1,89,1,4,
/* out0136_em-eta16-phi6*/	4,36,1,4,92,0,6,88,1,1,88,2,4,
/* out0137_em-eta17-phi6*/	7,36,0,1,36,1,3,92,0,2,105,1,3,88,0,2,88,1,1,88,2,2,
/* out0138_em-eta18-phi6*/	3,36,0,1,105,1,4,88,0,4,
/* out0139_em-eta19-phi6*/	2,105,0,2,105,1,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	1,116,3,14,
/* out0142_em-eta2-phi7*/	2,116,2,16,116,3,2,
/* out0143_em-eta3-phi7*/	2,115,2,2,115,3,16,
/* out0144_em-eta4-phi7*/	2,66,1,3,115,2,14,
/* out0145_em-eta5-phi7*/	8,64,0,3,64,1,1,64,2,14,65,0,5,65,1,2,66,0,16,66,1,9,66,2,2,
/* out0146_em-eta6-phi7*/	6,67,2,8,59,1,1,59,2,3,62,2,3,64,0,10,64,1,9,
/* out0147_em-eta7-phi7*/	7,67,0,9,67,1,10,67,2,6,58,2,3,59,1,7,62,0,12,62,2,1,
/* out0148_em-eta8-phi7*/	9,45,1,4,45,2,1,65,0,8,65,2,5,67,0,1,67,1,1,58,0,1,58,1,8,58,2,9,
/* out0149_em-eta9-phi7*/	8,44,1,1,44,2,9,45,1,1,65,0,7,57,0,1,57,2,7,58,0,1,58,1,7,
/* out0150_em-eta10-phi7*/	5,44,1,13,44,2,1,57,0,11,57,1,1,57,2,1,
/* out0151_em-eta11-phi7*/	11,43,0,2,43,2,9,44,1,1,95,0,10,95,1,1,95,2,5,56,0,1,57,0,3,57,1,1,90,1,2,90,2,4,
/* out0152_em-eta12-phi7*/	6,43,0,8,43,1,2,93,2,5,95,2,10,56,0,2,90,1,6,
/* out0153_em-eta13-phi7*/	11,37,1,2,37,2,2,42,0,1,42,2,1,43,0,1,43,1,1,93,0,5,93,1,1,93,2,5,89,2,7,90,1,1,
/* out0154_em-eta14-phi7*/	8,37,1,4,42,0,3,93,0,6,93,1,2,106,2,1,89,0,2,89,1,2,89,2,2,
/* out0155_em-eta15-phi7*/	9,36,1,3,36,2,2,42,0,1,92,0,2,92,2,1,106,1,4,106,2,1,89,0,2,89,1,4,
/* out0156_em-eta16-phi7*/	7,36,1,4,92,0,3,105,1,1,105,2,1,106,1,3,88,2,4,89,1,1,
/* out0157_em-eta17-phi7*/	5,36,0,5,36,1,1,105,1,4,105,2,1,88,2,4,
/* out0158_em-eta18-phi7*/	4,105,0,2,105,1,3,88,0,3,88,2,1,
/* out0159_em-eta19-phi7*/	1,105,0,4,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	1,118,0,14,
/* out0162_em-eta2-phi8*/	2,118,0,2,118,1,16,
/* out0163_em-eta3-phi8*/	2,117,0,16,117,1,2,
/* out0164_em-eta4-phi8*/	3,66,1,3,66,2,3,117,1,14,
/* out0165_em-eta5-phi8*/	6,60,0,2,60,1,7,60,2,14,64,0,1,66,1,1,66,2,11,
/* out0166_em-eta6-phi8*/	8,46,0,8,46,2,1,67,2,1,59,0,3,59,2,12,60,0,2,60,1,9,64,0,2,
/* out0167_em-eta7-phi8*/	9,45,2,5,46,0,3,46,2,14,67,0,6,58,2,1,59,0,11,59,1,8,59,2,1,92,2,2,
/* out0168_em-eta8-phi8*/	7,45,0,5,45,1,6,45,2,9,58,0,10,58,2,3,92,1,6,92,2,1,
/* out0169_em-eta9-phi8*/	8,39,1,1,44,0,3,44,2,6,45,0,2,45,1,5,58,0,4,91,1,3,91,2,9,
/* out0170_em-eta10-phi8*/	5,38,2,1,44,0,12,57,0,1,90,2,1,91,1,10,
/* out0171_em-eta11-phi8*/	10,38,1,5,38,2,4,43,0,2,44,0,1,44,1,1,95,0,6,95,1,8,108,1,2,90,0,1,90,2,10,
/* out0172_em-eta12-phi8*/	8,37,2,3,38,1,4,43,0,3,95,1,7,95,2,1,107,2,5,90,0,4,90,1,5,
/* out0173_em-eta13-phi8*/	9,37,1,1,37,2,7,93,0,3,107,1,7,107,2,1,89,0,1,89,2,3,90,0,1,90,1,2,
/* out0174_em-eta14-phi8*/	6,37,0,1,37,1,6,93,0,2,106,2,6,107,1,1,89,0,6,
/* out0175_em-eta15-phi8*/	7,36,2,4,37,1,3,106,0,1,106,1,3,106,2,4,49,2,1,89,0,4,
/* out0176_em-eta16-phi8*/	5,36,0,1,36,2,5,106,1,6,49,1,2,49,2,3,
/* out0177_em-eta17-phi8*/	3,36,0,6,105,2,6,49,1,4,
/* out0178_em-eta18-phi8*/	3,105,0,4,105,2,3,49,1,2,
/* out0179_em-eta19-phi8*/	1,105,0,3,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	1,118,3,14,
/* out0182_em-eta2-phi9*/	2,118,2,16,118,3,2,
/* out0183_em-eta3-phi9*/	2,117,2,2,117,3,16,
/* out0184_em-eta4-phi9*/	2,94,2,2,117,2,14,
/* out0185_em-eta5-phi9*/	4,60,0,8,60,2,2,94,1,11,94,2,7,
/* out0186_em-eta6-phi9*/	9,41,0,1,41,1,5,46,0,5,46,1,4,60,0,4,93,0,2,93,1,7,93,2,14,94,1,1,
/* out0187_em-eta7-phi9*/	9,40,2,9,41,1,2,45,2,1,46,1,12,46,2,1,59,0,2,92,0,1,92,2,11,93,1,9,
/* out0188_em-eta8-phi9*/	6,39,2,2,40,1,11,45,0,8,92,0,7,92,1,9,92,2,2,
/* out0189_em-eta9-phi9*/	8,39,0,1,39,1,5,39,2,11,45,0,1,52,1,1,91,0,6,91,2,7,92,1,1,
/* out0190_em-eta10-phi9*/	5,38,2,5,39,1,9,51,2,2,91,0,9,91,1,3,
/* out0191_em-eta11-phi9*/	9,38,0,4,38,1,2,38,2,6,108,0,6,108,1,10,51,1,4,51,2,1,90,0,4,90,2,1,
/* out0192_em-eta12-phi9*/	9,37,2,1,38,0,3,38,1,5,107,0,1,107,2,9,108,1,4,50,2,2,51,1,1,90,0,6,
/* out0193_em-eta13-phi9*/	7,37,0,5,37,2,3,107,0,5,107,1,5,107,2,1,50,1,2,50,2,5,
/* out0194_em-eta14-phi9*/	8,37,0,7,90,1,1,106,0,1,106,2,3,107,0,1,107,1,3,50,1,6,89,0,1,
/* out0195_em-eta15-phi9*/	8,31,1,1,31,2,2,36,2,1,37,0,1,106,0,7,106,2,1,49,2,4,50,1,1,
/* out0196_em-eta16-phi9*/	5,31,1,2,36,2,3,89,2,1,106,0,5,49,2,4,
/* out0197_em-eta17-phi9*/	7,31,1,1,36,0,2,36,2,1,89,1,2,89,2,1,105,2,2,49,1,4,
/* out0198_em-eta18-phi9*/	3,89,1,2,105,2,3,49,1,3,
/* out0199_em-eta19-phi9*/	1,105,0,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	1,120,0,14,
/* out0202_em-eta2-phi10*/	2,120,0,2,120,1,16,
/* out0203_em-eta3-phi10*/	2,119,0,16,119,1,2,
/* out0204_em-eta4-phi10*/	4,55,0,1,55,1,1,94,2,3,119,1,14,
/* out0205_em-eta5-phi10*/	5,54,2,5,55,1,7,94,0,16,94,1,3,94,2,4,
/* out0206_em-eta6-phi10*/	8,41,0,10,41,1,2,53,2,1,54,1,9,54,2,3,93,0,10,93,2,2,94,1,1,
/* out0207_em-eta7-phi10*/	10,35,1,3,35,2,2,40,0,5,40,2,7,41,0,4,41,1,7,53,1,7,53,2,10,92,0,2,93,0,4,
/* out0208_em-eta8-phi10*/	7,34,2,4,39,2,1,40,0,11,40,1,5,52,2,8,53,1,5,92,0,6,
/* out0209_em-eta9-phi10*/	5,34,1,5,39,0,10,39,2,2,52,1,10,52,2,5,
/* out0210_em-eta10-phi10*/	8,33,1,2,33,2,6,38,0,1,39,0,5,39,1,1,51,2,9,52,1,3,91,0,1,
/* out0211_em-eta11-phi10*/	7,33,1,5,38,0,6,91,2,3,108,0,9,51,0,2,51,1,6,51,2,3,
/* out0212_em-eta12-phi10*/	8,32,2,8,38,0,2,91,1,5,91,2,4,107,0,3,108,0,1,50,2,4,51,1,5,
/* out0213_em-eta13-phi10*/	8,32,1,8,37,0,1,90,2,3,91,1,2,107,0,6,50,0,3,50,1,1,50,2,4,
/* out0214_em-eta14-phi10*/	7,31,2,4,32,1,2,37,0,1,90,1,3,90,2,6,50,0,2,50,1,4,
/* out0215_em-eta15-phi10*/	7,31,1,1,31,2,5,90,1,6,106,0,1,49,0,1,49,2,3,50,1,2,
/* out0216_em-eta16-phi10*/	5,31,1,5,89,2,6,106,0,1,49,0,3,49,2,1,
/* out0217_em-eta17-phi10*/	4,31,1,2,89,1,3,89,2,3,49,0,3,
/* out0218_em-eta18-phi10*/	3,89,1,5,49,0,2,49,1,1,
/* out0219_em-eta19-phi10*/	1,89,1,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	1,120,3,14,
/* out0222_em-eta2-phi11*/	2,120,2,16,120,3,2,
/* out0223_em-eta3-phi11*/	2,119,2,2,119,3,16,
/* out0224_em-eta4-phi11*/	2,55,0,2,119,2,14,
/* out0225_em-eta5-phi11*/	5,48,0,7,54,0,3,54,2,6,55,0,13,55,1,8,
/* out0226_em-eta6-phi11*/	8,35,0,1,35,2,6,41,0,1,47,0,4,53,2,1,54,0,13,54,1,7,54,2,2,
/* out0227_em-eta7-phi11*/	7,35,0,8,35,1,9,35,2,8,47,0,3,53,0,13,53,1,1,53,2,4,
/* out0228_em-eta8-phi11*/	8,34,0,4,34,2,12,35,1,4,46,0,6,52,0,3,52,2,3,53,0,3,53,1,3,
/* out0229_em-eta9-phi11*/	7,33,2,1,34,0,5,34,1,11,45,0,1,46,0,1,52,0,12,52,1,1,
/* out0230_em-eta10-phi11*/	8,33,0,5,33,1,1,33,2,9,45,0,6,51,0,3,51,2,1,52,0,1,52,1,1,
/* out0231_em-eta11-phi11*/	7,32,2,1,33,0,3,33,1,8,91,0,1,91,2,6,44,0,1,51,0,9,
/* out0232_em-eta12-phi11*/	9,32,0,3,32,2,7,91,0,6,91,1,4,91,2,3,44,0,5,50,0,1,50,2,1,51,0,2,
/* out0233_em-eta13-phi11*/	8,32,0,5,32,1,3,90,0,1,90,2,4,91,0,1,91,1,5,44,0,2,50,0,6,
/* out0234_em-eta14-phi11*/	9,31,0,1,31,2,3,32,0,1,32,1,3,90,0,5,90,1,1,90,2,3,43,0,2,50,0,4,
/* out0235_em-eta15-phi11*/	6,31,0,4,31,2,2,90,0,3,90,1,5,43,0,4,49,0,1,
/* out0236_em-eta16-phi11*/	6,31,0,3,31,1,2,89,0,2,89,2,4,43,0,2,49,0,3,
/* out0237_em-eta17-phi11*/	6,31,0,1,31,1,2,89,0,4,89,2,1,42,0,1,49,0,3,
/* out0238_em-eta18-phi11*/	3,89,0,2,89,1,2,42,0,3,
/* out0239_em-eta19-phi11*/	2,89,1,1,42,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	1,122,0,14,
/* out0242_em-eta2-phi12*/	2,122,0,2,122,1,16,
/* out0243_em-eta3-phi12*/	2,121,0,16,121,1,2,
/* out0244_em-eta4-phi12*/	3,41,0,1,48,1,1,121,1,14,
/* out0245_em-eta5-phi12*/	4,41,0,2,48,0,8,48,1,14,48,2,10,
/* out0246_em-eta6-phi12*/	7,30,0,8,40,0,1,47,0,5,47,1,14,47,2,1,48,0,1,48,2,5,
/* out0247_em-eta7-phi12*/	9,29,0,4,29,1,5,30,0,6,30,2,6,35,0,7,46,0,1,46,1,6,47,0,4,47,2,12,
/* out0248_em-eta8-phi12*/	6,29,0,12,29,2,4,34,0,3,46,0,7,46,1,6,46,2,6,
/* out0249_em-eta9-phi12*/	7,28,0,9,28,1,3,34,0,4,45,0,2,45,1,8,46,0,1,46,2,5,
/* out0250_em-eta10-phi12*/	7,27,1,1,28,0,7,28,2,2,33,0,5,45,0,6,45,1,2,45,2,5,
/* out0251_em-eta11-phi12*/	9,27,0,8,27,1,1,33,0,3,88,0,9,91,0,1,44,0,1,44,1,5,45,0,1,45,2,4,
/* out0252_em-eta12-phi12*/	10,27,0,6,32,0,3,87,0,2,87,1,1,88,0,3,88,2,2,91,0,6,44,0,5,44,1,2,44,2,1,
/* out0253_em-eta13-phi12*/	8,26,0,3,26,1,1,32,0,4,87,0,9,91,0,1,43,1,1,44,0,2,44,2,5,
/* out0254_em-eta14-phi12*/	6,26,0,6,87,0,3,87,2,1,90,0,5,43,0,2,43,1,4,
/* out0255_em-eta15-phi12*/	6,26,0,2,31,0,4,86,0,5,90,0,2,43,0,4,43,2,1,
/* out0256_em-eta16-phi12*/	6,25,0,2,31,0,3,86,0,5,89,0,2,43,0,2,43,2,3,
/* out0257_em-eta17-phi12*/	5,25,0,2,25,1,1,86,0,1,89,0,4,42,0,4,
/* out0258_em-eta18-phi12*/	4,85,0,3,89,0,2,42,0,3,42,1,1,
/* out0259_em-eta19-phi12*/	2,85,1,1,42,1,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	1,122,3,14,
/* out0262_em-eta2-phi13*/	2,122,2,16,122,3,2,
/* out0263_em-eta3-phi13*/	2,121,2,2,121,3,16,
/* out0264_em-eta4-phi13*/	3,41,0,5,41,2,1,121,2,14,
/* out0265_em-eta5-phi13*/	6,40,0,4,40,1,11,41,0,8,41,2,13,48,1,1,48,2,1,
/* out0266_em-eta6-phi13*/	10,24,0,2,24,1,2,30,0,2,30,2,4,39,1,3,40,0,11,40,1,1,40,2,10,47,1,2,47,2,1,
/* out0267_em-eta7-phi13*/	8,24,0,12,29,1,8,30,2,6,39,0,14,39,1,4,39,2,2,46,1,1,47,2,2,
/* out0268_em-eta8-phi13*/	9,23,0,5,29,1,3,29,2,12,38,0,4,38,1,3,39,0,2,39,2,3,46,1,3,46,2,4,
/* out0269_em-eta9-phi13*/	6,23,0,2,28,1,12,28,2,2,38,0,11,45,1,3,46,2,1,
/* out0270_em-eta10-phi13*/	7,22,0,1,27,1,2,28,2,11,37,0,3,38,2,1,45,1,3,45,2,6,
/* out0271_em-eta11-phi13*/	8,27,0,1,27,1,9,27,2,1,88,0,4,88,2,7,37,0,5,44,1,4,45,2,1,
/* out0272_em-eta12-phi13*/	7,27,0,1,27,2,9,84,0,1,87,1,8,88,2,6,44,1,5,44,2,4,
/* out0273_em-eta13-phi13*/	9,26,0,1,26,1,7,27,2,1,87,0,2,87,1,4,87,2,5,36,0,2,43,1,1,44,2,5,
/* out0274_em-eta14-phi13*/	6,26,0,3,26,1,1,26,2,2,86,1,3,87,2,6,43,1,6,
/* out0275_em-eta15-phi13*/	7,25,0,1,26,0,1,26,2,4,86,0,2,86,1,5,43,1,2,43,2,4,
/* out0276_em-eta16-phi13*/	4,25,0,7,86,0,3,86,2,4,43,2,4,
/* out0277_em-eta17-phi13*/	6,25,0,1,25,1,2,85,0,4,86,2,2,42,0,4,42,1,1,
/* out0278_em-eta18-phi13*/	4,85,0,5,85,1,2,42,0,1,42,1,3,
/* out0279_em-eta19-phi13*/	1,85,1,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	1,124,0,14,
/* out0282_em-eta2-phi14*/	2,124,0,2,124,1,16,
/* out0283_em-eta3-phi14*/	2,123,0,16,123,1,2,
/* out0284_em-eta4-phi14*/	4,24,0,4,24,2,1,41,2,1,123,1,14,
/* out0285_em-eta5-phi14*/	6,23,1,1,24,0,9,24,1,10,24,2,15,40,1,3,41,2,1,
/* out0286_em-eta6-phi14*/	7,24,1,9,23,0,14,23,1,4,23,2,1,39,1,2,40,1,1,40,2,6,
/* out0287_em-eta7-phi14*/	11,18,0,3,23,1,1,24,0,2,24,1,5,24,2,16,22,0,4,22,1,1,23,0,2,23,2,1,39,1,7,39,2,8,
/* out0288_em-eta8-phi14*/	6,23,0,5,23,1,13,23,2,3,22,0,5,38,1,11,39,2,3,
/* out0289_em-eta9-phi14*/	9,22,0,1,22,1,4,23,0,4,23,2,8,28,1,1,28,2,1,38,0,1,38,1,2,38,2,13,
/* out0290_em-eta10-phi14*/	6,22,0,11,22,1,3,22,2,1,37,0,2,37,1,10,38,2,1,
/* out0291_em-eta11-phi14*/	12,21,0,1,21,1,1,22,0,3,22,2,2,27,1,3,27,2,2,84,0,5,84,1,7,88,2,1,37,0,5,37,1,1,37,2,5,
/* out0292_em-eta12-phi14*/	10,21,0,6,27,2,3,84,0,10,84,2,2,87,1,1,36,0,2,36,1,4,37,0,1,37,2,2,44,2,1,
/* out0293_em-eta13-phi14*/	8,21,0,3,26,1,6,82,0,3,82,1,1,84,2,1,87,1,2,87,2,3,36,0,7,
/* out0294_em-eta14-phi14*/	7,26,1,1,26,2,5,82,0,6,86,1,2,87,2,1,36,0,4,43,1,1,
/* out0295_em-eta15-phi14*/	10,20,0,1,25,0,1,25,1,1,26,2,4,82,0,1,86,1,6,86,2,2,35,0,2,43,1,1,43,2,3,
/* out0296_em-eta16-phi14*/	5,25,0,2,25,1,5,86,2,6,35,0,3,43,2,1,
/* out0297_em-eta17-phi14*/	6,25,1,2,85,0,3,85,1,2,86,2,1,35,0,1,42,1,3,
/* out0298_em-eta18-phi14*/	3,85,0,1,85,1,5,42,1,4,
/* out0299_em-eta19-phi14*/	0,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	1,124,3,14,
/* out0302_em-eta2-phi15*/	2,124,2,16,124,3,2,
/* out0303_em-eta3-phi15*/	2,123,2,2,123,3,16,
/* out0304_em-eta4-phi15*/	1,123,2,14,
/* out0305_em-eta5-phi15*/	6,23,1,2,24,0,3,24,1,6,28,0,14,28,1,7,28,2,1,
/* out0306_em-eta6-phi15*/	9,18,1,1,19,0,1,19,1,7,23,1,9,23,2,10,26,0,4,26,1,1,28,0,2,28,2,1,
/* out0307_em-eta7-phi15*/	8,18,0,9,18,1,12,18,2,4,22,0,2,22,1,14,22,2,1,23,2,4,26,0,2,
/* out0308_em-eta8-phi15*/	9,16,0,3,16,1,4,18,0,4,18,2,5,23,1,2,23,2,3,21,1,2,22,0,5,22,2,10,
/* out0309_em-eta9-phi15*/	6,16,0,11,22,1,4,23,2,2,21,0,10,21,1,4,38,2,1,
/* out0310_em-eta10-phi15*/	6,22,1,5,22,2,8,21,0,6,21,2,1,37,1,5,37,2,1,
/* out0311_em-eta11-phi15*/	7,15,0,1,21,1,6,22,2,5,84,1,9,84,2,1,20,0,4,37,2,7,
/* out0312_em-eta12-phi15*/	8,21,0,3,21,1,5,21,2,2,83,1,1,84,2,11,20,0,1,36,1,7,37,2,1,
/* out0313_em-eta13-phi15*/	9,20,1,1,21,0,3,21,2,5,82,0,1,82,1,10,84,2,1,36,0,1,36,1,3,36,2,4,
/* out0314_em-eta14-phi15*/	8,20,0,4,20,1,2,26,2,1,82,0,4,82,1,1,82,2,4,35,1,1,36,2,6,
/* out0315_em-eta15-phi15*/	8,20,0,6,81,0,1,81,1,2,82,0,1,82,2,3,86,2,1,35,0,1,35,1,4,
/* out0316_em-eta16-phi15*/	4,20,0,2,25,1,4,81,0,6,35,0,4,
/* out0317_em-eta17-phi15*/	4,25,1,1,81,0,5,85,1,1,35,0,4,
/* out0318_em-eta18-phi15*/	3,85,1,4,35,0,1,42,1,2,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	1,126,0,14,
/* out0322_em-eta2-phi16*/	2,126,0,2,126,1,16,
/* out0323_em-eta3-phi16*/	2,125,0,16,125,1,2,
/* out0324_em-eta4-phi16*/	2,28,1,1,125,1,14,
/* out0325_em-eta5-phi16*/	4,27,1,7,27,2,2,28,1,8,28,2,11,
/* out0326_em-eta6-phi16*/	8,19,0,4,19,1,9,19,2,12,26,0,4,26,1,14,26,2,4,27,1,3,28,2,3,
/* out0327_em-eta7-phi16*/	11,17,1,6,17,2,4,18,1,3,18,2,5,19,0,10,22,1,1,22,2,2,25,0,2,25,1,5,26,0,6,26,2,8,
/* out0328_em-eta8-phi16*/	7,16,1,11,16,2,1,17,1,7,18,2,2,21,1,3,22,2,3,25,0,12,
/* out0329_em-eta9-phi16*/	7,15,1,1,16,0,2,16,1,1,16,2,13,21,1,7,21,2,8,25,0,1,
/* out0330_em-eta10-phi16*/	5,15,0,6,15,1,7,16,2,1,20,1,6,21,2,7,
/* out0331_em-eta11-phi16*/	8,15,0,9,15,2,2,21,1,2,83,1,1,83,2,6,20,0,6,20,1,4,20,2,1,
/* out0332_em-eta12-phi16*/	9,11,1,1,21,1,2,21,2,5,83,0,1,83,1,10,83,2,2,20,0,5,20,2,2,36,1,2,
/* out0333_em-eta13-phi16*/	9,11,1,1,20,1,3,21,2,4,82,1,4,82,2,1,83,0,1,83,1,4,14,1,3,36,2,4,
/* out0334_em-eta14-phi16*/	6,20,1,7,79,0,2,82,2,7,14,1,2,35,1,2,36,2,2,
/* out0335_em-eta15-phi16*/	6,20,0,2,20,2,3,79,0,1,81,1,6,82,2,1,35,1,5,
/* out0336_em-eta16-phi16*/	7,20,0,1,20,2,3,81,0,1,81,1,4,81,2,1,35,1,1,35,2,3,
/* out0337_em-eta17-phi16*/	3,81,0,2,81,2,4,35,2,4,
/* out0338_em-eta18-phi16*/	3,81,0,1,81,2,1,35,2,1,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	1,126,3,14,
/* out0342_em-eta2-phi17*/	2,126,2,16,126,3,2,
/* out0343_em-eta3-phi17*/	2,125,2,2,125,3,16,
/* out0344_em-eta4-phi17*/	1,125,2,14,
/* out0345_em-eta5-phi17*/	3,27,0,9,27,1,3,27,2,14,
/* out0346_em-eta6-phi17*/	8,19,2,4,71,0,11,26,1,1,26,2,2,27,0,7,27,1,3,33,0,5,33,1,8,
/* out0347_em-eta7-phi17*/	10,17,0,6,17,1,1,17,2,12,19,0,1,71,1,1,71,2,16,25,1,9,25,2,1,26,2,2,33,0,10,
/* out0348_em-eta8-phi17*/	8,17,0,10,17,1,2,68,1,1,68,2,6,25,0,1,25,1,2,25,2,14,29,2,1,
/* out0349_em-eta9-phi17*/	7,15,1,1,16,2,1,68,1,13,68,2,1,25,2,1,29,1,7,29,2,7,
/* out0350_em-eta10-phi17*/	5,15,1,7,15,2,5,68,1,2,20,1,3,29,1,9,
/* out0351_em-eta11-phi17*/	5,11,2,2,15,2,9,83,2,5,20,1,3,20,2,8,
/* out0352_em-eta12-phi17*/	6,11,1,5,11,2,6,83,0,10,83,2,3,14,2,4,20,2,5,
/* out0353_em-eta13-phi17*/	5,11,1,8,79,1,6,83,0,4,14,1,4,14,2,4,
/* out0354_em-eta14-phi17*/	6,11,1,1,20,1,3,20,2,2,79,0,8,79,1,1,14,1,6,
/* out0355_em-eta15-phi17*/	6,20,2,6,79,0,5,81,1,3,14,1,1,35,1,3,35,2,1,
/* out0356_em-eta16-phi17*/	4,20,2,2,81,1,1,81,2,5,35,2,4,
/* out0357_em-eta17-phi17*/	2,81,2,5,35,2,3,
/* out0358_em-eta18-phi17*/	0,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	1,128,0,14,
/* out0362_em-eta2-phi18*/	2,128,0,2,128,1,16,
/* out0363_em-eta3-phi18*/	2,127,0,16,127,1,2,
/* out0364_em-eta4-phi18*/	1,127,1,14,
/* out0365_em-eta5-phi18*/	3,34,0,9,34,1,14,34,2,3,
/* out0366_em-eta6-phi18*/	10,70,1,10,70,2,1,71,0,5,71,1,7,31,1,2,31,2,1,33,1,8,33,2,5,34,0,7,34,2,3,
/* out0367_em-eta7-phi18*/	11,69,0,1,69,1,6,69,2,12,70,0,1,70,1,1,71,1,8,30,1,1,30,2,9,31,1,2,33,0,1,33,2,11,
/* out0368_em-eta8-phi18*/	8,68,0,1,68,2,7,69,0,2,69,1,10,29,2,1,30,0,1,30,1,14,30,2,2,
/* out0369_em-eta9-phi18*/	7,12,2,1,13,1,1,68,0,13,68,2,2,29,0,7,29,2,7,30,1,1,
/* out0370_em-eta10-phi18*/	5,12,1,5,12,2,7,68,0,2,15,2,3,29,0,9,
/* out0371_em-eta11-phi18*/	5,11,2,2,12,1,9,80,1,5,15,1,8,15,2,3,
/* out0372_em-eta12-phi18*/	6,11,0,4,11,2,6,80,0,10,80,1,3,14,2,4,15,1,5,
/* out0373_em-eta13-phi18*/	5,11,0,7,79,1,7,80,0,4,14,0,4,14,2,4,
/* out0374_em-eta14-phi18*/	6,6,1,2,6,2,3,11,0,1,79,1,2,79,2,7,14,0,6,
/* out0375_em-eta15-phi18*/	6,6,1,6,76,2,3,79,2,5,7,1,1,7,2,3,14,0,1,
/* out0376_em-eta16-phi18*/	4,6,1,2,76,1,5,76,2,1,7,1,4,
/* out0377_em-eta17-phi18*/	2,76,1,5,7,1,3,
/* out0378_em-eta18-phi18*/	0,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	1,128,3,14,
/* out0382_em-eta2-phi19*/	2,128,2,16,128,3,2,
/* out0383_em-eta3-phi19*/	2,127,2,2,127,3,16,
/* out0384_em-eta4-phi19*/	2,32,2,1,127,2,14,
/* out0385_em-eta5-phi19*/	4,32,1,11,32,2,8,34,1,2,34,2,7,
/* out0386_em-eta6-phi19*/	8,70,0,4,70,1,5,70,2,13,31,0,4,31,1,4,31,2,14,32,1,3,34,2,3,
/* out0387_em-eta7-phi19*/	11,14,1,5,14,2,3,69,0,6,69,2,4,70,0,10,17,1,2,17,2,1,30,0,2,30,2,5,31,0,6,31,1,8,
/* out0388_em-eta8-phi19*/	7,13,1,1,13,2,11,14,1,2,69,0,7,16,2,3,17,1,3,30,0,12,
/* out0389_em-eta9-phi19*/	7,12,2,1,13,0,2,13,1,13,13,2,1,16,1,8,16,2,7,30,0,1,
/* out0390_em-eta10-phi19*/	5,12,0,6,12,2,7,13,1,1,15,2,6,16,1,7,
/* out0391_em-eta11-phi19*/	8,7,2,2,12,0,9,12,1,2,80,1,6,80,2,1,15,0,6,15,1,1,15,2,4,
/* out0392_em-eta12-phi19*/	9,7,1,5,7,2,2,11,0,2,80,0,1,80,1,2,80,2,10,8,2,2,15,0,5,15,1,2,
/* out0393_em-eta13-phi19*/	10,6,2,3,7,1,4,11,0,2,77,1,1,77,2,4,79,2,1,80,0,1,80,2,4,8,1,4,14,0,3,
/* out0394_em-eta14-phi19*/	6,6,2,7,77,1,7,79,2,2,7,2,2,8,1,2,14,0,2,
/* out0395_em-eta15-phi19*/	6,6,0,2,6,1,3,76,2,6,77,1,1,79,2,1,7,2,5,
/* out0396_em-eta16-phi19*/	7,6,0,1,6,1,3,76,0,1,76,1,1,76,2,4,7,1,3,7,2,1,
/* out0397_em-eta17-phi19*/	3,76,0,2,76,1,4,7,1,4,
/* out0398_em-eta18-phi19*/	3,76,0,1,76,1,1,7,1,1,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	1,130,0,14,
/* out0402_em-eta2-phi20*/	2,130,0,2,130,1,16,
/* out0403_em-eta3-phi20*/	2,129,0,16,129,1,2,
/* out0404_em-eta4-phi20*/	1,129,1,14,
/* out0405_em-eta5-phi20*/	6,18,2,2,19,0,3,19,2,7,32,0,14,32,1,1,32,2,7,
/* out0406_em-eta6-phi20*/	9,14,2,1,70,0,1,70,2,2,18,1,10,18,2,9,31,0,4,31,2,1,32,0,2,32,1,1,
/* out0407_em-eta7-phi20*/	8,14,0,9,14,1,4,14,2,12,17,0,2,17,1,1,17,2,14,18,1,4,31,0,2,
/* out0408_em-eta8-phi20*/	9,9,1,3,9,2,2,13,0,3,13,2,4,14,0,4,14,1,5,16,2,2,17,0,5,17,1,10,
/* out0409_em-eta9-phi20*/	6,8,2,4,9,1,2,13,0,11,10,1,1,16,0,10,16,2,4,
/* out0410_em-eta10-phi20*/	6,8,1,8,8,2,5,9,1,1,9,2,5,16,0,6,16,1,1,
/* out0411_em-eta11-phi20*/	7,7,2,6,8,1,5,12,0,1,78,1,1,78,2,9,9,1,7,15,0,4,
/* out0412_em-eta12-phi20*/	8,7,0,3,7,1,2,7,2,5,78,1,11,80,2,1,8,2,7,9,1,1,15,0,1,
/* out0413_em-eta13-phi20*/	9,6,2,1,7,0,3,7,1,5,77,0,1,77,2,10,78,1,1,8,0,1,8,1,4,8,2,3,
/* out0414_em-eta14-phi20*/	8,1,1,1,6,0,4,6,2,2,77,0,4,77,1,4,77,2,1,7,2,1,8,1,6,
/* out0415_em-eta15-phi20*/	8,6,0,6,73,1,1,76,0,1,76,2,2,77,0,1,77,1,3,7,0,1,7,2,4,
/* out0416_em-eta16-phi20*/	4,0,1,4,6,0,2,76,0,6,7,0,4,
/* out0417_em-eta17-phi20*/	4,0,1,1,72,1,1,76,0,5,7,0,4,
/* out0418_em-eta18-phi20*/	3,72,1,4,0,1,2,7,0,1,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	1,130,3,14,
/* out0422_em-eta2-phi21*/	2,130,2,16,130,3,2,
/* out0423_em-eta3-phi21*/	2,129,2,2,129,3,16,
/* out0424_em-eta4-phi21*/	4,13,1,1,19,0,4,19,1,1,129,2,14,
/* out0425_em-eta5-phi21*/	6,12,2,3,13,1,1,18,2,1,19,0,9,19,1,15,19,2,9,
/* out0426_em-eta6-phi21*/	7,10,2,9,11,2,2,12,1,6,12,2,1,18,0,14,18,1,1,18,2,4,
/* out0427_em-eta7-phi21*/	11,9,2,1,10,0,2,10,1,16,10,2,5,14,0,3,11,1,8,11,2,7,17,0,4,17,2,1,18,0,2,18,1,1,
/* out0428_em-eta8-phi21*/	6,9,0,5,9,1,3,9,2,13,10,2,11,11,1,3,17,0,5,
/* out0429_em-eta9-phi21*/	9,3,1,1,3,2,1,8,0,1,8,2,4,9,0,4,9,1,8,10,0,1,10,1,13,10,2,2,
/* out0430_em-eta10-phi21*/	6,8,0,11,8,1,1,8,2,3,9,0,2,9,2,10,10,1,1,
/* out0431_em-eta11-phi21*/	12,2,1,2,2,2,3,7,0,1,7,2,1,8,0,3,8,1,2,75,1,1,78,0,5,78,2,7,9,0,5,9,1,5,9,2,1,
/* out0432_em-eta12-phi21*/	10,2,1,3,7,0,6,74,2,1,78,0,10,78,1,2,2,1,1,8,0,2,8,2,4,9,0,1,9,1,2,
/* out0433_em-eta13-phi21*/	8,1,2,6,7,0,3,74,1,3,74,2,2,77,0,3,77,2,1,78,1,1,8,0,7,
/* out0434_em-eta14-phi21*/	7,1,1,5,1,2,1,73,2,2,74,1,1,77,0,6,1,2,1,8,0,4,
/* out0435_em-eta15-phi21*/	10,0,1,1,0,2,1,1,1,4,6,0,1,73,1,2,73,2,6,77,0,1,1,1,3,1,2,1,7,0,2,
/* out0436_em-eta16-phi21*/	6,0,1,5,0,2,2,73,1,6,0,2,1,1,1,1,7,0,3,
/* out0437_em-eta17-phi21*/	7,0,1,2,72,1,2,72,2,3,73,1,1,0,1,3,0,2,1,7,0,1,
/* out0438_em-eta18-phi21*/	3,72,1,5,72,2,1,0,1,4,
/* out0439_em-eta19-phi21*/	0,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	1,132,0,14,
/* out0442_em-eta2-phi22*/	2,132,0,2,132,1,16,
/* out0443_em-eta3-phi22*/	2,131,0,16,131,1,2,
/* out0444_em-eta4-phi22*/	3,13,0,5,13,1,1,131,1,14,
/* out0445_em-eta5-phi22*/	6,6,1,1,6,2,1,12,0,4,12,2,11,13,0,8,13,1,13,
/* out0446_em-eta6-phi22*/	10,5,0,2,5,1,4,10,0,2,10,2,2,5,1,1,5,2,2,11,2,3,12,0,11,12,1,10,12,2,1,
/* out0447_em-eta7-phi22*/	8,4,2,8,5,1,6,10,0,12,4,2,1,5,1,2,11,0,14,11,1,2,11,2,4,
/* out0448_em-eta8-phi22*/	9,4,1,12,4,2,3,9,0,5,4,1,4,4,2,3,10,0,4,10,2,3,11,0,2,11,1,3,
/* out0449_em-eta9-phi22*/	6,3,1,2,3,2,12,9,0,2,3,2,3,4,1,1,10,0,11,
/* out0450_em-eta10-phi22*/	7,2,2,2,3,1,11,8,0,1,3,1,6,3,2,3,9,0,3,10,1,1,
/* out0451_em-eta11-phi22*/	8,2,0,1,2,1,1,2,2,9,75,0,4,75,1,7,2,2,4,3,1,1,9,0,5,
/* out0452_em-eta12-phi22*/	7,2,0,1,2,1,9,74,2,8,75,1,6,78,0,1,2,1,4,2,2,5,
/* out0453_em-eta13-phi22*/	9,1,0,1,1,2,7,2,1,1,74,0,2,74,1,5,74,2,4,1,2,1,2,1,5,8,0,2,
/* out0454_em-eta14-phi22*/	6,1,0,3,1,1,2,1,2,1,73,2,3,74,1,6,1,2,6,
/* out0455_em-eta15-phi22*/	7,0,2,1,1,0,1,1,1,4,73,0,2,73,2,5,1,1,4,1,2,2,
/* out0456_em-eta16-phi22*/	5,0,2,7,73,0,3,73,1,4,0,2,1,1,1,4,
/* out0457_em-eta17-phi22*/	6,0,1,2,0,2,1,72,2,4,73,1,2,0,1,1,0,2,4,
/* out0458_em-eta18-phi22*/	4,72,1,2,72,2,5,0,1,4,0,2,1,
/* out0459_em-eta19-phi22*/	1,72,1,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	1,132,3,14,
/* out0462_em-eta2-phi23*/	2,132,2,16,132,3,2,
/* out0463_em-eta3-phi23*/	2,131,2,2,131,3,16,
/* out0464_em-eta4-phi23*/	4,6,0,7,6,2,1,13,0,1,131,2,14,
/* out0465_em-eta5-phi23*/	4,6,0,8,6,1,10,6,2,14,13,0,2,
/* out0466_em-eta6-phi23*/	7,5,0,8,5,0,5,5,1,1,5,2,14,6,0,1,6,1,5,12,0,1,
/* out0467_em-eta7-phi23*/	8,4,0,4,4,2,5,5,0,6,5,1,6,4,0,8,4,2,6,5,0,11,5,1,12,
/* out0468_em-eta8-phi23*/	5,4,0,12,4,1,4,4,0,7,4,1,6,4,2,6,
/* out0469_em-eta9-phi23*/	6,3,0,9,3,2,3,3,0,2,3,2,8,4,0,1,4,1,5,
/* out0470_em-eta10-phi23*/	6,2,2,1,3,0,7,3,1,2,3,0,13,3,1,5,3,2,2,
/* out0471_em-eta11-phi23*/	7,2,0,8,2,2,1,75,0,9,2,0,8,2,2,5,3,0,1,3,1,4,
/* out0472_em-eta12-phi23*/	8,2,0,6,74,0,2,74,2,1,75,0,3,75,1,2,2,0,6,2,1,1,2,2,2,
/* out0473_em-eta13-phi23*/	7,1,0,3,1,2,1,74,0,9,1,0,5,1,2,1,2,0,2,2,1,5,
/* out0474_em-eta14-phi23*/	5,1,0,6,74,0,3,74,1,1,1,0,3,1,2,4,
/* out0475_em-eta15-phi23*/	4,1,0,2,73,0,5,1,0,5,1,1,1,
/* out0476_em-eta16-phi23*/	4,0,2,2,73,0,5,1,0,2,1,1,3,
/* out0477_em-eta17-phi23*/	5,0,1,1,0,2,2,73,0,1,0,2,5,1,0,1,
/* out0478_em-eta18-phi23*/	3,72,2,3,0,1,1,0,2,3,
/* out0479_em-eta19-phi23*/	2,72,1,1,0,1,1
};