parameter integer matrixH [0:4944] = {
/* num inputs = 155(in0-in154) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 8 */
//* total number of input in adders 1488 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	1, 99, 0, 13, 
/* out0002_had-eta2-phi0*/	2, 99, 0, 3, 99, 1, 14, 
/* out0003_had-eta3-phi0*/	2, 98, 0, 16, 99, 1, 2, 
/* out0004_had-eta4-phi0*/	3, 87, 0, 1, 87, 1, 1, 98, 1, 16, 
/* out0005_had-eta5-phi0*/	5, 86, 2, 10, 87, 0, 2, 87, 1, 14, 97, 0, 16, 97, 1, 2, 
/* out0006_had-eta6-phi0*/	6, 85, 2, 1, 86, 0, 1, 86, 1, 14, 86, 2, 5, 96, 0, 2, 97, 1, 14, 
/* out0007_had-eta7-phi0*/	4, 85, 1, 6, 85, 2, 12, 96, 0, 14, 96, 1, 4, 
/* out0008_had-eta8-phi0*/	4, 84, 2, 6, 85, 1, 6, 96, 1, 12, 96, 2, 4, 
/* out0009_had-eta9-phi0*/	4, 84, 1, 8, 84, 2, 5, 95, 0, 3, 96, 2, 12, 
/* out0010_had-eta10-phi0*/	4, 83, 2, 5, 84, 1, 2, 95, 0, 13, 95, 1, 3, 
/* out0011_had-eta11-phi0*/	3, 83, 1, 5, 83, 2, 4, 95, 1, 13, 
/* out0012_had-eta12-phi0*/	2, 82, 2, 1, 83, 1, 2, 
/* out0013_had-eta13-phi0*/	2, 82, 1, 1, 82, 2, 5, 
/* out0014_had-eta14-phi0*/	1, 82, 1, 4, 
/* out0015_had-eta15-phi0*/	1, 81, 2, 1, 
/* out0016_had-eta16-phi0*/	1, 81, 2, 3, 
/* out0017_had-eta17-phi0*/	1, 81, 1, 2, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	1, 99, 3, 13, 
/* out0022_had-eta2-phi1*/	2, 99, 2, 14, 99, 3, 3, 
/* out0023_had-eta3-phi1*/	2, 98, 3, 16, 99, 2, 2, 
/* out0024_had-eta4-phi1*/	3, 80, 2, 3, 87, 0, 3, 98, 2, 16, 
/* out0025_had-eta5-phi1*/	8, 80, 1, 11, 80, 2, 11, 86, 0, 4, 86, 2, 1, 87, 0, 10, 87, 1, 1, 97, 2, 2, 97, 3, 16, 
/* out0026_had-eta6-phi1*/	8, 79, 1, 3, 79, 2, 10, 80, 1, 1, 85, 2, 1, 86, 0, 11, 86, 1, 2, 96, 5, 2, 97, 2, 14, 
/* out0027_had-eta7-phi1*/	7, 78, 2, 2, 79, 1, 4, 85, 0, 14, 85, 1, 1, 85, 2, 2, 96, 4, 4, 96, 5, 14, 
/* out0028_had-eta8-phi1*/	8, 78, 1, 3, 78, 2, 3, 84, 0, 4, 84, 2, 4, 85, 0, 2, 85, 1, 3, 96, 3, 4, 96, 4, 12, 
/* out0029_had-eta9-phi1*/	5, 84, 0, 11, 84, 1, 3, 84, 2, 1, 95, 3, 3, 96, 3, 12, 
/* out0030_had-eta10-phi1*/	6, 77, 2, 1, 83, 0, 3, 83, 2, 6, 84, 1, 3, 95, 2, 3, 95, 3, 13, 
/* out0031_had-eta11-phi1*/	4, 83, 0, 5, 83, 1, 4, 83, 2, 1, 95, 2, 13, 
/* out0032_had-eta12-phi1*/	2, 82, 2, 4, 83, 1, 5, 
/* out0033_had-eta13-phi1*/	3, 82, 0, 2, 82, 1, 1, 82, 2, 5, 
/* out0034_had-eta14-phi1*/	1, 82, 1, 6, 
/* out0035_had-eta15-phi1*/	2, 81, 2, 4, 82, 1, 2, 
/* out0036_had-eta16-phi1*/	1, 81, 2, 4, 
/* out0037_had-eta17-phi1*/	1, 81, 1, 4, 
/* out0038_had-eta18-phi1*/	1, 81, 1, 3, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	1, 104, 0, 13, 
/* out0042_had-eta2-phi2*/	2, 104, 0, 3, 104, 1, 14, 
/* out0043_had-eta3-phi2*/	2, 103, 0, 16, 104, 1, 2, 
/* out0044_had-eta4-phi2*/	3, 80, 0, 1, 80, 2, 1, 103, 1, 16, 
/* out0045_had-eta5-phi2*/	7, 74, 1, 1, 74, 2, 9, 80, 0, 15, 80, 1, 3, 80, 2, 1, 102, 0, 16, 102, 1, 2, 
/* out0046_had-eta6-phi2*/	8, 73, 2, 1, 74, 1, 4, 79, 0, 14, 79, 1, 2, 79, 2, 6, 80, 1, 1, 101, 0, 2, 102, 1, 14, 
/* out0047_had-eta7-phi2*/	8, 73, 1, 1, 73, 2, 1, 78, 0, 4, 78, 2, 8, 79, 0, 2, 79, 1, 7, 101, 0, 14, 101, 1, 4, 
/* out0048_had-eta8-phi2*/	5, 78, 0, 4, 78, 1, 11, 78, 2, 3, 101, 1, 12, 101, 2, 4, 
/* out0049_had-eta9-phi2*/	5, 77, 2, 13, 78, 1, 2, 84, 0, 1, 100, 0, 3, 101, 2, 12, 
/* out0050_had-eta10-phi2*/	5, 77, 1, 10, 77, 2, 1, 83, 0, 2, 100, 0, 13, 100, 1, 3, 
/* out0051_had-eta11-phi2*/	4, 76, 2, 5, 77, 1, 1, 83, 0, 5, 100, 1, 13, 
/* out0052_had-eta12-phi2*/	5, 76, 1, 4, 76, 2, 2, 82, 0, 2, 82, 2, 1, 83, 0, 1, 
/* out0053_had-eta13-phi2*/	1, 82, 0, 7, 
/* out0054_had-eta14-phi2*/	2, 82, 0, 4, 82, 1, 1, 
/* out0055_had-eta15-phi2*/	3, 81, 0, 2, 81, 2, 3, 82, 1, 1, 
/* out0056_had-eta16-phi2*/	2, 81, 0, 3, 81, 2, 1, 
/* out0057_had-eta17-phi2*/	2, 81, 0, 1, 81, 1, 3, 
/* out0058_had-eta18-phi2*/	1, 81, 1, 3, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 104, 3, 13, 
/* out0062_had-eta2-phi3*/	2, 104, 2, 14, 104, 3, 3, 
/* out0063_had-eta3-phi3*/	2, 103, 3, 16, 104, 2, 2, 
/* out0064_had-eta4-phi3*/	2, 69, 2, 14, 103, 2, 16, 
/* out0065_had-eta5-phi3*/	8, 68, 2, 1, 69, 1, 7, 69, 2, 2, 74, 0, 14, 74, 1, 2, 74, 2, 7, 102, 2, 2, 102, 3, 16, 
/* out0066_had-eta6-phi3*/	8, 68, 1, 1, 68, 2, 1, 73, 0, 4, 73, 2, 10, 74, 0, 2, 74, 1, 9, 101, 5, 2, 102, 2, 14, 
/* out0067_had-eta7-phi3*/	7, 72, 2, 1, 73, 0, 2, 73, 1, 14, 73, 2, 4, 78, 0, 2, 101, 4, 4, 101, 5, 14, 
/* out0068_had-eta8-phi3*/	5, 72, 1, 2, 72, 2, 10, 78, 0, 6, 101, 3, 4, 101, 4, 12, 
/* out0069_had-eta9-phi3*/	5, 72, 1, 4, 77, 0, 10, 77, 2, 1, 100, 3, 3, 101, 3, 12, 
/* out0070_had-eta10-phi3*/	6, 71, 2, 1, 76, 2, 1, 77, 0, 6, 77, 1, 5, 100, 2, 3, 100, 3, 13, 
/* out0071_had-eta11-phi3*/	3, 76, 0, 4, 76, 2, 7, 100, 2, 13, 
/* out0072_had-eta12-phi3*/	3, 76, 0, 1, 76, 1, 7, 76, 2, 1, 
/* out0073_had-eta13-phi3*/	3, 75, 2, 4, 76, 1, 3, 82, 0, 1, 
/* out0074_had-eta14-phi3*/	2, 75, 1, 1, 75, 2, 6, 
/* out0075_had-eta15-phi3*/	2, 75, 1, 4, 81, 0, 1, 
/* out0076_had-eta16-phi3*/	1, 81, 0, 4, 
/* out0077_had-eta17-phi3*/	1, 81, 0, 4, 
/* out0078_had-eta18-phi3*/	2, 81, 0, 1, 81, 1, 1, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 109, 0, 13, 
/* out0082_had-eta2-phi4*/	2, 109, 0, 3, 109, 1, 14, 
/* out0083_had-eta3-phi4*/	2, 108, 0, 16, 109, 1, 2, 
/* out0084_had-eta4-phi4*/	4, 69, 0, 6, 69, 1, 1, 70, 2, 1, 108, 1, 16, 
/* out0085_had-eta5-phi4*/	8, 68, 0, 7, 68, 2, 11, 69, 0, 10, 69, 1, 8, 70, 1, 2, 70, 2, 11, 107, 0, 16, 107, 1, 2, 
/* out0086_had-eta6-phi4*/	7, 67, 2, 4, 68, 0, 3, 68, 1, 14, 68, 2, 3, 73, 0, 4, 106, 0, 2, 107, 1, 14, 
/* out0087_had-eta7-phi4*/	8, 67, 1, 5, 67, 2, 8, 72, 0, 2, 72, 2, 2, 73, 0, 6, 73, 1, 1, 106, 0, 14, 106, 1, 4, 
/* out0088_had-eta8-phi4*/	5, 72, 0, 12, 72, 1, 3, 72, 2, 3, 106, 1, 12, 106, 2, 4, 
/* out0089_had-eta9-phi4*/	5, 71, 2, 8, 72, 0, 1, 72, 1, 7, 105, 0, 3, 106, 2, 12, 
/* out0090_had-eta10-phi4*/	4, 71, 1, 6, 71, 2, 7, 105, 0, 13, 105, 1, 3, 
/* out0091_had-eta11-phi4*/	4, 56, 2, 1, 71, 1, 3, 76, 0, 6, 105, 1, 13, 
/* out0092_had-eta12-phi4*/	3, 56, 2, 2, 76, 0, 5, 76, 1, 2, 
/* out0093_had-eta13-phi4*/	2, 75, 0, 3, 75, 2, 4, 
/* out0094_had-eta14-phi4*/	3, 75, 0, 2, 75, 1, 2, 75, 2, 2, 
/* out0095_had-eta15-phi4*/	1, 75, 1, 5, 
/* out0096_had-eta16-phi4*/	2, 75, 1, 1, 88, 2, 3, 
/* out0097_had-eta17-phi4*/	1, 88, 2, 3, 
/* out0098_had-eta18-phi4*/	2, 88, 1, 2, 88, 2, 1, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 109, 3, 13, 
/* out0102_had-eta2-phi5*/	2, 109, 2, 14, 109, 3, 3, 
/* out0103_had-eta3-phi5*/	2, 108, 3, 16, 109, 2, 2, 
/* out0104_had-eta4-phi5*/	1, 108, 2, 16, 
/* out0105_had-eta5-phi5*/	7, 63, 2, 9, 68, 0, 3, 70, 0, 16, 70, 1, 14, 70, 2, 4, 107, 2, 2, 107, 3, 16, 
/* out0106_had-eta6-phi5*/	8, 63, 1, 8, 63, 2, 7, 67, 0, 5, 67, 2, 2, 68, 0, 3, 68, 1, 1, 106, 5, 2, 107, 2, 14, 
/* out0107_had-eta7-phi5*/	6, 61, 2, 1, 67, 0, 11, 67, 1, 9, 67, 2, 2, 106, 4, 4, 106, 5, 14, 
/* out0108_had-eta8-phi5*/	6, 61, 1, 1, 61, 2, 14, 67, 1, 2, 72, 0, 1, 106, 3, 4, 106, 4, 12, 
/* out0109_had-eta9-phi5*/	5, 61, 1, 7, 61, 2, 1, 71, 0, 7, 105, 3, 3, 106, 3, 12, 
/* out0110_had-eta10-phi5*/	4, 71, 0, 9, 71, 1, 4, 105, 2, 3, 105, 3, 13, 
/* out0111_had-eta11-phi5*/	3, 56, 2, 8, 71, 1, 3, 105, 2, 13, 
/* out0112_had-eta12-phi5*/	2, 56, 1, 4, 56, 2, 5, 
/* out0113_had-eta13-phi5*/	2, 56, 1, 4, 75, 0, 4, 
/* out0114_had-eta14-phi5*/	1, 75, 0, 6, 
/* out0115_had-eta15-phi5*/	3, 75, 0, 1, 75, 1, 3, 88, 2, 1, 
/* out0116_had-eta16-phi5*/	1, 88, 2, 5, 
/* out0117_had-eta17-phi5*/	2, 88, 1, 1, 88, 2, 3, 
/* out0118_had-eta18-phi5*/	1, 88, 1, 5, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 114, 0, 13, 
/* out0122_had-eta2-phi6*/	2, 114, 0, 3, 114, 1, 14, 
/* out0123_had-eta3-phi6*/	2, 113, 0, 16, 114, 1, 2, 
/* out0124_had-eta4-phi6*/	1, 113, 1, 16, 
/* out0125_had-eta5-phi6*/	7, 63, 0, 9, 64, 2, 3, 65, 0, 4, 65, 1, 14, 65, 2, 16, 112, 0, 16, 112, 1, 2, 
/* out0126_had-eta6-phi6*/	8, 62, 0, 2, 62, 2, 5, 63, 0, 7, 63, 1, 8, 64, 1, 1, 64, 2, 3, 111, 0, 2, 112, 1, 14, 
/* out0127_had-eta7-phi6*/	6, 61, 0, 1, 62, 0, 2, 62, 1, 9, 62, 2, 11, 111, 0, 14, 111, 1, 4, 
/* out0128_had-eta8-phi6*/	6, 58, 2, 1, 61, 0, 14, 61, 1, 1, 62, 1, 2, 111, 1, 12, 111, 2, 4, 
/* out0129_had-eta9-phi6*/	5, 57, 2, 7, 61, 0, 1, 61, 1, 7, 110, 0, 3, 111, 2, 12, 
/* out0130_had-eta10-phi6*/	4, 57, 1, 4, 57, 2, 9, 110, 0, 13, 110, 1, 3, 
/* out0131_had-eta11-phi6*/	3, 56, 0, 8, 57, 1, 3, 110, 1, 13, 
/* out0132_had-eta12-phi6*/	2, 56, 0, 5, 56, 1, 4, 
/* out0133_had-eta13-phi6*/	2, 56, 1, 4, 89, 2, 4, 
/* out0134_had-eta14-phi6*/	1, 89, 2, 6, 
/* out0135_had-eta15-phi6*/	3, 88, 0, 1, 89, 1, 3, 89, 2, 1, 
/* out0136_had-eta16-phi6*/	1, 88, 0, 4, 
/* out0137_had-eta17-phi6*/	2, 88, 0, 3, 88, 1, 1, 
/* out0138_had-eta18-phi6*/	1, 88, 1, 5, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 114, 3, 13, 
/* out0142_had-eta2-phi7*/	2, 114, 2, 14, 114, 3, 3, 
/* out0143_had-eta3-phi7*/	2, 113, 3, 16, 114, 2, 2, 
/* out0144_had-eta4-phi7*/	4, 65, 0, 1, 66, 1, 1, 66, 2, 6, 113, 2, 16, 
/* out0145_had-eta5-phi7*/	8, 64, 0, 11, 64, 2, 7, 65, 0, 11, 65, 1, 2, 66, 1, 8, 66, 2, 10, 112, 2, 2, 112, 3, 16, 
/* out0146_had-eta6-phi7*/	7, 59, 2, 4, 62, 0, 4, 64, 0, 3, 64, 1, 14, 64, 2, 3, 111, 5, 2, 112, 2, 14, 
/* out0147_had-eta7-phi7*/	8, 58, 0, 2, 58, 2, 2, 59, 1, 1, 59, 2, 6, 62, 0, 8, 62, 1, 5, 111, 4, 4, 111, 5, 14, 
/* out0148_had-eta8-phi7*/	5, 58, 0, 3, 58, 1, 3, 58, 2, 12, 111, 3, 4, 111, 4, 12, 
/* out0149_had-eta9-phi7*/	5, 57, 0, 8, 58, 1, 7, 58, 2, 1, 110, 3, 3, 111, 3, 12, 
/* out0150_had-eta10-phi7*/	4, 57, 0, 7, 57, 1, 6, 110, 2, 3, 110, 3, 13, 
/* out0151_had-eta11-phi7*/	4, 56, 0, 1, 57, 1, 3, 90, 2, 6, 110, 2, 13, 
/* out0152_had-eta12-phi7*/	3, 56, 0, 2, 90, 1, 2, 90, 2, 5, 
/* out0153_had-eta13-phi7*/	2, 89, 0, 4, 89, 2, 3, 
/* out0154_had-eta14-phi7*/	3, 89, 0, 2, 89, 1, 2, 89, 2, 2, 
/* out0155_had-eta15-phi7*/	1, 89, 1, 5, 
/* out0156_had-eta16-phi7*/	2, 88, 0, 3, 89, 1, 1, 
/* out0157_had-eta17-phi7*/	1, 88, 0, 4, 
/* out0158_had-eta18-phi7*/	2, 88, 0, 1, 88, 1, 2, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 119, 0, 13, 
/* out0162_had-eta2-phi8*/	2, 119, 0, 3, 119, 1, 14, 
/* out0163_had-eta3-phi8*/	2, 118, 0, 16, 119, 1, 2, 
/* out0164_had-eta4-phi8*/	2, 66, 0, 14, 118, 1, 16, 
/* out0165_had-eta5-phi8*/	8, 60, 0, 7, 60, 1, 2, 60, 2, 14, 64, 0, 1, 66, 0, 2, 66, 1, 7, 117, 0, 16, 117, 1, 2, 
/* out0166_had-eta6-phi8*/	8, 59, 0, 10, 59, 2, 4, 60, 1, 9, 60, 2, 2, 64, 0, 1, 64, 1, 1, 116, 0, 2, 117, 1, 14, 
/* out0167_had-eta7-phi8*/	7, 58, 0, 1, 59, 0, 4, 59, 1, 14, 59, 2, 2, 92, 2, 2, 116, 0, 14, 116, 1, 4, 
/* out0168_had-eta8-phi8*/	5, 58, 0, 10, 58, 1, 2, 92, 2, 6, 116, 1, 12, 116, 2, 4, 
/* out0169_had-eta9-phi8*/	5, 58, 1, 4, 91, 0, 1, 91, 2, 10, 115, 0, 3, 116, 2, 12, 
/* out0170_had-eta10-phi8*/	6, 57, 0, 1, 90, 0, 1, 91, 1, 5, 91, 2, 6, 115, 0, 13, 115, 1, 3, 
/* out0171_had-eta11-phi8*/	3, 90, 0, 7, 90, 2, 4, 115, 1, 13, 
/* out0172_had-eta12-phi8*/	3, 90, 0, 1, 90, 1, 7, 90, 2, 1, 
/* out0173_had-eta13-phi8*/	3, 50, 2, 1, 89, 0, 4, 90, 1, 3, 
/* out0174_had-eta14-phi8*/	2, 89, 0, 6, 89, 1, 1, 
/* out0175_had-eta15-phi8*/	2, 49, 2, 1, 89, 1, 4, 
/* out0176_had-eta16-phi8*/	1, 49, 2, 4, 
/* out0177_had-eta17-phi8*/	1, 49, 2, 4, 
/* out0178_had-eta18-phi8*/	2, 49, 1, 1, 49, 2, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 119, 3, 13, 
/* out0182_had-eta2-phi9*/	2, 119, 2, 14, 119, 3, 3, 
/* out0183_had-eta3-phi9*/	2, 118, 3, 16, 119, 2, 2, 
/* out0184_had-eta4-phi9*/	3, 94, 0, 1, 94, 2, 1, 118, 2, 16, 
/* out0185_had-eta5-phi9*/	7, 60, 0, 9, 60, 1, 1, 94, 0, 1, 94, 1, 3, 94, 2, 15, 117, 2, 2, 117, 3, 16, 
/* out0186_had-eta6-phi9*/	8, 59, 0, 1, 60, 1, 4, 93, 0, 6, 93, 1, 2, 93, 2, 14, 94, 1, 1, 116, 5, 2, 117, 2, 14, 
/* out0187_had-eta7-phi9*/	8, 59, 0, 1, 59, 1, 1, 92, 0, 8, 92, 2, 4, 93, 1, 7, 93, 2, 2, 116, 4, 4, 116, 5, 14, 
/* out0188_had-eta8-phi9*/	5, 92, 0, 3, 92, 1, 11, 92, 2, 4, 116, 3, 4, 116, 4, 12, 
/* out0189_had-eta9-phi9*/	5, 52, 2, 1, 91, 0, 13, 92, 1, 2, 115, 3, 3, 116, 3, 12, 
/* out0190_had-eta10-phi9*/	5, 51, 2, 2, 91, 0, 1, 91, 1, 10, 115, 2, 3, 115, 3, 13, 
/* out0191_had-eta11-phi9*/	4, 51, 2, 5, 90, 0, 5, 91, 1, 1, 115, 2, 13, 
/* out0192_had-eta12-phi9*/	5, 50, 0, 1, 50, 2, 2, 51, 2, 1, 90, 0, 2, 90, 1, 4, 
/* out0193_had-eta13-phi9*/	1, 50, 2, 7, 
/* out0194_had-eta14-phi9*/	2, 50, 1, 1, 50, 2, 4, 
/* out0195_had-eta15-phi9*/	3, 49, 0, 3, 49, 2, 2, 50, 1, 1, 
/* out0196_had-eta16-phi9*/	2, 49, 0, 1, 49, 2, 3, 
/* out0197_had-eta17-phi9*/	2, 49, 1, 3, 49, 2, 1, 
/* out0198_had-eta18-phi9*/	1, 49, 1, 3, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 124, 0, 13, 
/* out0202_had-eta2-phi10*/	2, 124, 0, 3, 124, 1, 14, 
/* out0203_had-eta3-phi10*/	2, 123, 0, 16, 124, 1, 2, 
/* out0204_had-eta4-phi10*/	3, 55, 1, 3, 94, 0, 3, 123, 1, 16, 
/* out0205_had-eta5-phi10*/	8, 54, 0, 1, 54, 2, 4, 55, 0, 1, 55, 1, 10, 94, 0, 11, 94, 1, 11, 122, 0, 16, 122, 1, 2, 
/* out0206_had-eta6-phi10*/	8, 53, 0, 1, 54, 1, 2, 54, 2, 11, 93, 0, 10, 93, 1, 3, 94, 1, 1, 121, 0, 2, 122, 1, 14, 
/* out0207_had-eta7-phi10*/	7, 53, 0, 2, 53, 1, 1, 53, 2, 14, 92, 0, 2, 93, 1, 4, 121, 0, 14, 121, 1, 4, 
/* out0208_had-eta8-phi10*/	8, 52, 0, 4, 52, 2, 4, 53, 1, 3, 53, 2, 2, 92, 0, 3, 92, 1, 3, 121, 1, 12, 121, 2, 4, 
/* out0209_had-eta9-phi10*/	5, 52, 0, 1, 52, 1, 3, 52, 2, 11, 120, 0, 3, 121, 2, 12, 
/* out0210_had-eta10-phi10*/	6, 51, 0, 6, 51, 2, 3, 52, 1, 3, 91, 0, 1, 120, 0, 13, 120, 1, 3, 
/* out0211_had-eta11-phi10*/	4, 51, 0, 1, 51, 1, 4, 51, 2, 5, 120, 1, 13, 
/* out0212_had-eta12-phi10*/	2, 50, 0, 4, 51, 1, 5, 
/* out0213_had-eta13-phi10*/	3, 50, 0, 5, 50, 1, 1, 50, 2, 2, 
/* out0214_had-eta14-phi10*/	1, 50, 1, 6, 
/* out0215_had-eta15-phi10*/	2, 49, 0, 4, 50, 1, 2, 
/* out0216_had-eta16-phi10*/	1, 49, 0, 4, 
/* out0217_had-eta17-phi10*/	1, 49, 1, 4, 
/* out0218_had-eta18-phi10*/	1, 49, 1, 3, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 124, 3, 13, 
/* out0222_had-eta2-phi11*/	2, 124, 2, 14, 124, 3, 3, 
/* out0223_had-eta3-phi11*/	2, 123, 3, 16, 124, 2, 2, 
/* out0224_had-eta4-phi11*/	3, 55, 0, 1, 55, 1, 1, 123, 2, 16, 
/* out0225_had-eta5-phi11*/	6, 48, 2, 7, 54, 0, 10, 55, 0, 14, 55, 1, 2, 122, 2, 2, 122, 3, 16, 
/* out0226_had-eta6-phi11*/	7, 47, 2, 4, 53, 0, 1, 54, 0, 5, 54, 1, 14, 54, 2, 1, 121, 5, 2, 122, 2, 14, 
/* out0227_had-eta7-phi11*/	5, 47, 2, 3, 53, 0, 12, 53, 1, 6, 121, 4, 4, 121, 5, 14, 
/* out0228_had-eta8-phi11*/	5, 46, 2, 6, 52, 0, 6, 53, 1, 6, 121, 3, 4, 121, 4, 12, 
/* out0229_had-eta9-phi11*/	6, 45, 2, 1, 46, 2, 1, 52, 0, 5, 52, 1, 8, 120, 3, 3, 121, 3, 12, 
/* out0230_had-eta10-phi11*/	5, 45, 2, 6, 51, 0, 5, 52, 1, 2, 120, 2, 3, 120, 3, 13, 
/* out0231_had-eta11-phi11*/	4, 44, 2, 1, 51, 0, 4, 51, 1, 5, 120, 2, 13, 
/* out0232_had-eta12-phi11*/	3, 44, 2, 5, 50, 0, 1, 51, 1, 2, 
/* out0233_had-eta13-phi11*/	3, 44, 2, 2, 50, 0, 5, 50, 1, 1, 
/* out0234_had-eta14-phi11*/	2, 43, 2, 2, 50, 1, 4, 
/* out0235_had-eta15-phi11*/	2, 43, 2, 4, 49, 0, 1, 
/* out0236_had-eta16-phi11*/	2, 43, 2, 2, 49, 0, 3, 
/* out0237_had-eta17-phi11*/	2, 42, 1, 2, 49, 1, 2, 
/* out0238_had-eta18-phi11*/	1, 42, 1, 5, 
/* out0239_had-eta19-phi11*/	1, 42, 1, 1, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 129, 0, 13, 
/* out0242_had-eta2-phi12*/	2, 129, 0, 3, 129, 1, 14, 
/* out0243_had-eta3-phi12*/	2, 128, 0, 16, 129, 1, 2, 
/* out0244_had-eta4-phi12*/	3, 41, 1, 1, 48, 0, 1, 128, 1, 16, 
/* out0245_had-eta5-phi12*/	6, 41, 1, 2, 48, 0, 14, 48, 1, 10, 48, 2, 8, 127, 0, 16, 127, 1, 2, 
/* out0246_had-eta6-phi12*/	8, 40, 2, 1, 47, 0, 14, 47, 1, 1, 47, 2, 5, 48, 1, 5, 48, 2, 1, 126, 0, 2, 127, 1, 14, 
/* out0247_had-eta7-phi12*/	6, 46, 0, 6, 46, 2, 1, 47, 1, 12, 47, 2, 4, 126, 0, 14, 126, 1, 4, 
/* out0248_had-eta8-phi12*/	5, 46, 0, 6, 46, 1, 6, 46, 2, 7, 126, 1, 12, 126, 2, 4, 
/* out0249_had-eta9-phi12*/	6, 45, 0, 8, 45, 2, 2, 46, 1, 5, 46, 2, 1, 125, 0, 3, 126, 2, 12, 
/* out0250_had-eta10-phi12*/	5, 45, 0, 2, 45, 1, 5, 45, 2, 6, 125, 0, 13, 125, 1, 3, 
/* out0251_had-eta11-phi12*/	5, 44, 0, 5, 44, 2, 1, 45, 1, 4, 45, 2, 1, 125, 1, 13, 
/* out0252_had-eta12-phi12*/	3, 44, 0, 2, 44, 1, 1, 44, 2, 5, 
/* out0253_had-eta13-phi12*/	3, 43, 0, 1, 44, 1, 5, 44, 2, 2, 
/* out0254_had-eta14-phi12*/	2, 43, 0, 4, 43, 2, 2, 
/* out0255_had-eta15-phi12*/	2, 43, 1, 1, 43, 2, 4, 
/* out0256_had-eta16-phi12*/	2, 43, 1, 3, 43, 2, 2, 
/* out0257_had-eta17-phi12*/	2, 42, 0, 2, 42, 1, 2, 
/* out0258_had-eta18-phi12*/	1, 42, 1, 5, 
/* out0259_had-eta19-phi12*/	1, 42, 1, 1, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 129, 3, 13, 
/* out0262_had-eta2-phi13*/	2, 129, 2, 14, 129, 3, 3, 
/* out0263_had-eta3-phi13*/	2, 128, 3, 16, 129, 2, 2, 
/* out0264_had-eta4-phi13*/	3, 41, 0, 3, 41, 1, 3, 128, 2, 16, 
/* out0265_had-eta5-phi13*/	8, 40, 0, 11, 40, 2, 4, 41, 0, 11, 41, 1, 10, 48, 0, 1, 48, 1, 1, 127, 2, 2, 127, 3, 16, 
/* out0266_had-eta6-phi13*/	8, 39, 0, 3, 40, 0, 1, 40, 1, 10, 40, 2, 11, 47, 0, 2, 47, 1, 1, 126, 5, 2, 127, 2, 14, 
/* out0267_had-eta7-phi13*/	7, 39, 0, 4, 39, 1, 2, 39, 2, 14, 46, 0, 1, 47, 1, 2, 126, 4, 4, 126, 5, 14, 
/* out0268_had-eta8-phi13*/	8, 38, 0, 3, 38, 2, 4, 39, 1, 3, 39, 2, 2, 46, 0, 3, 46, 1, 4, 126, 3, 4, 126, 4, 12, 
/* out0269_had-eta9-phi13*/	5, 38, 2, 11, 45, 0, 3, 46, 1, 1, 125, 3, 3, 126, 3, 12, 
/* out0270_had-eta10-phi13*/	6, 37, 2, 3, 38, 1, 1, 45, 0, 3, 45, 1, 6, 125, 2, 3, 125, 3, 13, 
/* out0271_had-eta11-phi13*/	4, 37, 2, 5, 44, 0, 4, 45, 1, 1, 125, 2, 13, 
/* out0272_had-eta12-phi13*/	2, 44, 0, 5, 44, 1, 4, 
/* out0273_had-eta13-phi13*/	3, 36, 2, 2, 43, 0, 1, 44, 1, 5, 
/* out0274_had-eta14-phi13*/	1, 43, 0, 6, 
/* out0275_had-eta15-phi13*/	2, 43, 0, 2, 43, 1, 4, 
/* out0276_had-eta16-phi13*/	1, 43, 1, 4, 
/* out0277_had-eta17-phi13*/	1, 42, 0, 4, 
/* out0278_had-eta18-phi13*/	1, 42, 0, 3, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 134, 0, 13, 
/* out0282_had-eta2-phi14*/	2, 134, 0, 3, 134, 1, 14, 
/* out0283_had-eta3-phi14*/	2, 133, 0, 16, 134, 1, 2, 
/* out0284_had-eta4-phi14*/	4, 24, 0, 4, 24, 2, 1, 41, 0, 1, 133, 1, 16, 
/* out0285_had-eta5-phi14*/	8, 23, 0, 1, 24, 0, 9, 24, 1, 9, 24, 2, 15, 40, 0, 3, 41, 0, 1, 132, 0, 16, 132, 1, 2, 
/* out0286_had-eta6-phi14*/	8, 23, 0, 4, 23, 1, 1, 23, 2, 14, 39, 0, 2, 40, 0, 1, 40, 1, 6, 131, 0, 2, 132, 1, 14, 
/* out0287_had-eta7-phi14*/	8, 22, 0, 1, 22, 2, 4, 23, 1, 1, 23, 2, 2, 39, 0, 7, 39, 1, 8, 131, 0, 14, 131, 1, 4, 
/* out0288_had-eta8-phi14*/	5, 22, 2, 5, 38, 0, 11, 39, 1, 3, 131, 1, 12, 131, 2, 4, 
/* out0289_had-eta9-phi14*/	5, 38, 0, 2, 38, 1, 13, 38, 2, 1, 130, 0, 3, 131, 2, 12, 
/* out0290_had-eta10-phi14*/	5, 37, 0, 10, 37, 2, 2, 38, 1, 1, 130, 0, 13, 130, 1, 3, 
/* out0291_had-eta11-phi14*/	4, 37, 0, 1, 37, 1, 5, 37, 2, 5, 130, 1, 13, 
/* out0292_had-eta12-phi14*/	5, 36, 0, 4, 36, 2, 2, 37, 1, 2, 37, 2, 1, 44, 1, 1, 
/* out0293_had-eta13-phi14*/	1, 36, 2, 7, 
/* out0294_had-eta14-phi14*/	2, 36, 2, 4, 43, 0, 1, 
/* out0295_had-eta15-phi14*/	3, 35, 2, 2, 43, 0, 1, 43, 1, 3, 
/* out0296_had-eta16-phi14*/	2, 35, 2, 3, 43, 1, 1, 
/* out0297_had-eta17-phi14*/	2, 35, 2, 1, 42, 0, 3, 
/* out0298_had-eta18-phi14*/	1, 42, 0, 3, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 134, 3, 13, 
/* out0302_had-eta2-phi15*/	2, 134, 2, 14, 134, 3, 3, 
/* out0303_had-eta3-phi15*/	2, 133, 3, 16, 134, 2, 2, 
/* out0304_had-eta4-phi15*/	1, 133, 2, 16, 
/* out0305_had-eta5-phi15*/	8, 23, 0, 2, 24, 0, 3, 24, 1, 7, 28, 0, 7, 28, 1, 1, 28, 2, 14, 132, 2, 2, 132, 3, 16, 
/* out0306_had-eta6-phi15*/	8, 23, 0, 9, 23, 1, 10, 26, 0, 1, 26, 2, 4, 28, 1, 1, 28, 2, 2, 131, 5, 2, 132, 2, 14, 
/* out0307_had-eta7-phi15*/	7, 22, 0, 14, 22, 1, 1, 22, 2, 2, 23, 1, 4, 26, 2, 2, 131, 4, 4, 131, 5, 14, 
/* out0308_had-eta8-phi15*/	5, 21, 0, 2, 22, 1, 10, 22, 2, 5, 131, 3, 4, 131, 4, 12, 
/* out0309_had-eta9-phi15*/	5, 21, 0, 4, 21, 2, 10, 38, 1, 1, 130, 3, 3, 131, 3, 12, 
/* out0310_had-eta10-phi15*/	6, 21, 1, 1, 21, 2, 6, 37, 0, 5, 37, 1, 1, 130, 2, 3, 130, 3, 13, 
/* out0311_had-eta11-phi15*/	3, 20, 2, 4, 37, 1, 7, 130, 2, 13, 
/* out0312_had-eta12-phi15*/	3, 20, 2, 1, 36, 0, 7, 37, 1, 1, 
/* out0313_had-eta13-phi15*/	3, 36, 0, 3, 36, 1, 4, 36, 2, 1, 
/* out0314_had-eta14-phi15*/	2, 35, 0, 1, 36, 1, 6, 
/* out0315_had-eta15-phi15*/	2, 35, 0, 4, 35, 2, 1, 
/* out0316_had-eta16-phi15*/	1, 35, 2, 4, 
/* out0317_had-eta17-phi15*/	1, 35, 2, 4, 
/* out0318_had-eta18-phi15*/	2, 35, 2, 1, 42, 0, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 139, 0, 13, 
/* out0322_had-eta2-phi16*/	2, 139, 0, 3, 139, 1, 14, 
/* out0323_had-eta3-phi16*/	2, 138, 0, 16, 139, 1, 2, 
/* out0324_had-eta4-phi16*/	2, 28, 0, 1, 138, 1, 16, 
/* out0325_had-eta5-phi16*/	6, 27, 0, 2, 27, 2, 7, 28, 0, 8, 28, 1, 11, 137, 0, 16, 137, 1, 2, 
/* out0326_had-eta6-phi16*/	7, 26, 0, 14, 26, 1, 4, 26, 2, 4, 27, 2, 3, 28, 1, 3, 136, 0, 2, 137, 1, 14, 
/* out0327_had-eta7-phi16*/	8, 22, 0, 1, 22, 1, 2, 25, 0, 5, 25, 2, 2, 26, 1, 8, 26, 2, 6, 136, 0, 14, 136, 1, 4, 
/* out0328_had-eta8-phi16*/	5, 21, 0, 3, 22, 1, 3, 25, 2, 12, 136, 1, 12, 136, 2, 4, 
/* out0329_had-eta9-phi16*/	5, 21, 0, 7, 21, 1, 8, 25, 2, 1, 135, 0, 3, 136, 2, 12, 
/* out0330_had-eta10-phi16*/	4, 20, 0, 6, 21, 1, 7, 135, 0, 13, 135, 1, 3, 
/* out0331_had-eta11-phi16*/	4, 20, 0, 4, 20, 1, 1, 20, 2, 6, 135, 1, 13, 
/* out0332_had-eta12-phi16*/	3, 20, 1, 2, 20, 2, 5, 36, 0, 2, 
/* out0333_had-eta13-phi16*/	2, 14, 2, 3, 36, 1, 4, 
/* out0334_had-eta14-phi16*/	3, 14, 2, 2, 35, 0, 2, 36, 1, 2, 
/* out0335_had-eta15-phi16*/	1, 35, 0, 5, 
/* out0336_had-eta16-phi16*/	2, 35, 0, 1, 35, 1, 3, 
/* out0337_had-eta17-phi16*/	1, 35, 1, 4, 
/* out0338_had-eta18-phi16*/	1, 35, 1, 1, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 139, 3, 13, 
/* out0342_had-eta2-phi17*/	2, 139, 2, 14, 139, 3, 3, 
/* out0343_had-eta3-phi17*/	2, 138, 3, 16, 139, 2, 2, 
/* out0344_had-eta4-phi17*/	1, 138, 2, 16, 
/* out0345_had-eta5-phi17*/	5, 27, 0, 14, 27, 1, 9, 27, 2, 3, 137, 2, 2, 137, 3, 16, 
/* out0346_had-eta6-phi17*/	8, 26, 0, 1, 26, 1, 2, 27, 1, 7, 27, 2, 3, 33, 0, 8, 33, 2, 5, 136, 5, 2, 137, 2, 14, 
/* out0347_had-eta7-phi17*/	6, 25, 0, 9, 25, 1, 1, 26, 1, 2, 33, 2, 10, 136, 4, 4, 136, 5, 14, 
/* out0348_had-eta8-phi17*/	6, 25, 0, 2, 25, 1, 14, 25, 2, 1, 29, 0, 1, 136, 3, 4, 136, 4, 12, 
/* out0349_had-eta9-phi17*/	5, 25, 1, 1, 29, 0, 7, 29, 2, 7, 135, 3, 3, 136, 3, 12, 
/* out0350_had-eta10-phi17*/	4, 20, 0, 3, 29, 2, 9, 135, 2, 3, 135, 3, 13, 
/* out0351_had-eta11-phi17*/	3, 20, 0, 3, 20, 1, 8, 135, 2, 13, 
/* out0352_had-eta12-phi17*/	2, 14, 0, 4, 20, 1, 5, 
/* out0353_had-eta13-phi17*/	2, 14, 0, 4, 14, 2, 4, 
/* out0354_had-eta14-phi17*/	1, 14, 2, 6, 
/* out0355_had-eta15-phi17*/	3, 14, 2, 1, 35, 0, 3, 35, 1, 1, 
/* out0356_had-eta16-phi17*/	1, 35, 1, 4, 
/* out0357_had-eta17-phi17*/	1, 35, 1, 3, 
/* out0358_had-eta18-phi17*/	0, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 144, 0, 13, 
/* out0362_had-eta2-phi18*/	2, 144, 0, 3, 144, 1, 14, 
/* out0363_had-eta3-phi18*/	2, 143, 0, 16, 144, 1, 2, 
/* out0364_had-eta4-phi18*/	1, 143, 1, 16, 
/* out0365_had-eta5-phi18*/	5, 34, 0, 14, 34, 1, 3, 34, 2, 9, 142, 0, 16, 142, 1, 2, 
/* out0366_had-eta6-phi18*/	8, 31, 0, 1, 31, 2, 2, 33, 0, 8, 33, 1, 5, 34, 1, 3, 34, 2, 7, 141, 0, 2, 142, 1, 14, 
/* out0367_had-eta7-phi18*/	7, 30, 0, 9, 30, 2, 1, 31, 2, 2, 33, 1, 11, 33, 2, 1, 141, 0, 14, 141, 1, 4, 
/* out0368_had-eta8-phi18*/	6, 29, 0, 1, 30, 0, 2, 30, 1, 1, 30, 2, 14, 141, 1, 12, 141, 2, 4, 
/* out0369_had-eta9-phi18*/	5, 29, 0, 7, 29, 1, 7, 30, 2, 1, 140, 0, 3, 141, 2, 12, 
/* out0370_had-eta10-phi18*/	4, 15, 0, 3, 29, 1, 9, 140, 0, 13, 140, 1, 3, 
/* out0371_had-eta11-phi18*/	3, 15, 0, 3, 15, 2, 8, 140, 1, 13, 
/* out0372_had-eta12-phi18*/	2, 14, 0, 4, 15, 2, 5, 
/* out0373_had-eta13-phi18*/	2, 14, 0, 4, 14, 1, 4, 
/* out0374_had-eta14-phi18*/	1, 14, 1, 6, 
/* out0375_had-eta15-phi18*/	3, 7, 0, 3, 7, 2, 1, 14, 1, 1, 
/* out0376_had-eta16-phi18*/	1, 7, 2, 4, 
/* out0377_had-eta17-phi18*/	1, 7, 2, 3, 
/* out0378_had-eta18-phi18*/	0, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 144, 3, 13, 
/* out0382_had-eta2-phi19*/	2, 144, 2, 14, 144, 3, 3, 
/* out0383_had-eta3-phi19*/	2, 143, 3, 16, 144, 2, 2, 
/* out0384_had-eta4-phi19*/	2, 32, 0, 1, 143, 2, 16, 
/* out0385_had-eta5-phi19*/	6, 32, 0, 8, 32, 2, 11, 34, 0, 2, 34, 1, 7, 142, 2, 2, 142, 3, 16, 
/* out0386_had-eta6-phi19*/	7, 31, 0, 14, 31, 1, 4, 31, 2, 4, 32, 2, 3, 34, 1, 3, 141, 5, 2, 142, 2, 14, 
/* out0387_had-eta7-phi19*/	8, 17, 0, 1, 17, 2, 2, 30, 0, 5, 30, 1, 2, 31, 1, 6, 31, 2, 8, 141, 4, 4, 141, 5, 14, 
/* out0388_had-eta8-phi19*/	5, 16, 0, 3, 17, 2, 3, 30, 1, 12, 141, 3, 4, 141, 4, 12, 
/* out0389_had-eta9-phi19*/	5, 16, 0, 7, 16, 2, 8, 30, 1, 1, 140, 3, 3, 141, 3, 12, 
/* out0390_had-eta10-phi19*/	4, 15, 0, 6, 16, 2, 7, 140, 2, 3, 140, 3, 13, 
/* out0391_had-eta11-phi19*/	4, 15, 0, 4, 15, 1, 6, 15, 2, 1, 140, 2, 13, 
/* out0392_had-eta12-phi19*/	3, 8, 0, 2, 15, 1, 5, 15, 2, 2, 
/* out0393_had-eta13-phi19*/	2, 8, 2, 4, 14, 1, 3, 
/* out0394_had-eta14-phi19*/	3, 7, 0, 2, 8, 2, 2, 14, 1, 2, 
/* out0395_had-eta15-phi19*/	1, 7, 0, 5, 
/* out0396_had-eta16-phi19*/	2, 7, 0, 1, 7, 2, 3, 
/* out0397_had-eta17-phi19*/	1, 7, 2, 4, 
/* out0398_had-eta18-phi19*/	1, 7, 2, 1, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 149, 0, 13, 
/* out0402_had-eta2-phi20*/	2, 149, 0, 3, 149, 1, 14, 
/* out0403_had-eta3-phi20*/	2, 148, 0, 16, 149, 1, 2, 
/* out0404_had-eta4-phi20*/	1, 148, 1, 16, 
/* out0405_had-eta5-phi20*/	8, 18, 0, 2, 19, 0, 3, 19, 2, 7, 32, 0, 7, 32, 1, 14, 32, 2, 1, 147, 0, 16, 147, 1, 2, 
/* out0406_had-eta6-phi20*/	8, 18, 0, 9, 18, 2, 10, 31, 0, 1, 31, 1, 4, 32, 1, 2, 32, 2, 1, 146, 0, 2, 147, 1, 14, 
/* out0407_had-eta7-phi20*/	7, 17, 0, 14, 17, 1, 2, 17, 2, 1, 18, 2, 4, 31, 1, 2, 146, 0, 14, 146, 1, 4, 
/* out0408_had-eta8-phi20*/	5, 16, 0, 2, 17, 1, 5, 17, 2, 10, 146, 1, 12, 146, 2, 4, 
/* out0409_had-eta9-phi20*/	5, 10, 2, 1, 16, 0, 4, 16, 1, 10, 145, 0, 3, 146, 2, 12, 
/* out0410_had-eta10-phi20*/	6, 9, 0, 5, 9, 2, 1, 16, 1, 6, 16, 2, 1, 145, 0, 13, 145, 1, 3, 
/* out0411_had-eta11-phi20*/	3, 9, 2, 7, 15, 1, 4, 145, 1, 13, 
/* out0412_had-eta12-phi20*/	3, 8, 0, 7, 9, 2, 1, 15, 1, 1, 
/* out0413_had-eta13-phi20*/	3, 8, 0, 3, 8, 1, 1, 8, 2, 4, 
/* out0414_had-eta14-phi20*/	2, 7, 0, 1, 8, 2, 6, 
/* out0415_had-eta15-phi20*/	2, 7, 0, 4, 7, 1, 1, 
/* out0416_had-eta16-phi20*/	1, 7, 1, 4, 
/* out0417_had-eta17-phi20*/	1, 7, 1, 4, 
/* out0418_had-eta18-phi20*/	2, 0, 0, 1, 7, 1, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 149, 3, 13, 
/* out0422_had-eta2-phi21*/	2, 149, 2, 14, 149, 3, 3, 
/* out0423_had-eta3-phi21*/	2, 148, 3, 16, 149, 2, 2, 
/* out0424_had-eta4-phi21*/	4, 13, 1, 1, 19, 0, 4, 19, 1, 1, 148, 2, 16, 
/* out0425_had-eta5-phi21*/	8, 12, 0, 3, 13, 1, 1, 18, 0, 1, 19, 0, 9, 19, 1, 15, 19, 2, 9, 147, 2, 2, 147, 3, 16, 
/* out0426_had-eta6-phi21*/	8, 11, 0, 2, 12, 0, 1, 12, 2, 6, 18, 0, 4, 18, 1, 14, 18, 2, 1, 146, 5, 2, 147, 2, 14, 
/* out0427_had-eta7-phi21*/	8, 11, 0, 7, 11, 2, 8, 17, 0, 1, 17, 1, 4, 18, 1, 2, 18, 2, 1, 146, 4, 4, 146, 5, 14, 
/* out0428_had-eta8-phi21*/	5, 10, 0, 11, 11, 2, 3, 17, 1, 5, 146, 3, 4, 146, 4, 12, 
/* out0429_had-eta9-phi21*/	5, 10, 0, 2, 10, 1, 1, 10, 2, 13, 145, 3, 3, 146, 3, 12, 
/* out0430_had-eta10-phi21*/	5, 9, 0, 10, 9, 1, 2, 10, 2, 1, 145, 2, 3, 145, 3, 13, 
/* out0431_had-eta11-phi21*/	4, 9, 0, 1, 9, 1, 5, 9, 2, 5, 145, 2, 13, 
/* out0432_had-eta12-phi21*/	5, 2, 2, 1, 8, 0, 4, 8, 1, 2, 9, 1, 1, 9, 2, 2, 
/* out0433_had-eta13-phi21*/	1, 8, 1, 7, 
/* out0434_had-eta14-phi21*/	2, 1, 0, 1, 8, 1, 4, 
/* out0435_had-eta15-phi21*/	3, 1, 0, 1, 1, 2, 3, 7, 1, 2, 
/* out0436_had-eta16-phi21*/	2, 1, 2, 1, 7, 1, 3, 
/* out0437_had-eta17-phi21*/	2, 0, 0, 3, 7, 1, 1, 
/* out0438_had-eta18-phi21*/	1, 0, 0, 3, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 154, 0, 13, 
/* out0442_had-eta2-phi22*/	2, 154, 0, 3, 154, 1, 14, 
/* out0443_had-eta3-phi22*/	2, 153, 0, 16, 154, 1, 2, 
/* out0444_had-eta4-phi22*/	3, 13, 0, 3, 13, 1, 3, 153, 1, 16, 
/* out0445_had-eta5-phi22*/	8, 6, 0, 1, 6, 2, 1, 12, 0, 11, 12, 1, 4, 13, 0, 10, 13, 1, 11, 152, 0, 16, 152, 1, 2, 
/* out0446_had-eta6-phi22*/	8, 5, 0, 2, 5, 2, 1, 11, 0, 3, 12, 0, 1, 12, 1, 11, 12, 2, 10, 151, 0, 2, 152, 1, 14, 
/* out0447_had-eta7-phi22*/	7, 4, 0, 1, 5, 2, 2, 11, 0, 4, 11, 1, 14, 11, 2, 2, 151, 0, 14, 151, 1, 4, 
/* out0448_had-eta8-phi22*/	8, 4, 0, 3, 4, 2, 4, 10, 0, 3, 10, 1, 4, 11, 1, 2, 11, 2, 3, 151, 1, 12, 151, 2, 4, 
/* out0449_had-eta9-phi22*/	5, 3, 0, 3, 4, 2, 1, 10, 1, 11, 150, 0, 3, 151, 2, 12, 
/* out0450_had-eta10-phi22*/	6, 3, 0, 3, 3, 2, 6, 9, 1, 3, 10, 2, 1, 150, 0, 13, 150, 1, 3, 
/* out0451_had-eta11-phi22*/	4, 2, 0, 4, 3, 2, 1, 9, 1, 5, 150, 1, 13, 
/* out0452_had-eta12-phi22*/	2, 2, 0, 5, 2, 2, 4, 
/* out0453_had-eta13-phi22*/	3, 1, 0, 1, 2, 2, 5, 8, 1, 2, 
/* out0454_had-eta14-phi22*/	1, 1, 0, 6, 
/* out0455_had-eta15-phi22*/	2, 1, 0, 2, 1, 2, 4, 
/* out0456_had-eta16-phi22*/	1, 1, 2, 4, 
/* out0457_had-eta17-phi22*/	1, 0, 0, 4, 
/* out0458_had-eta18-phi22*/	2, 0, 0, 3, 0, 1, 1, 
/* out0459_had-eta19-phi22*/	1, 0, 1, 6, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 154, 3, 13, 
/* out0462_had-eta2-phi23*/	2, 154, 2, 14, 154, 3, 3, 
/* out0463_had-eta3-phi23*/	2, 153, 3, 16, 154, 2, 2, 
/* out0464_had-eta4-phi23*/	4, 6, 0, 1, 6, 1, 7, 13, 0, 1, 153, 2, 16, 
/* out0465_had-eta5-phi23*/	6, 6, 0, 14, 6, 1, 8, 6, 2, 10, 13, 0, 2, 152, 2, 2, 152, 3, 16, 
/* out0466_had-eta6-phi23*/	8, 5, 0, 14, 5, 1, 5, 5, 2, 1, 6, 1, 1, 6, 2, 5, 12, 1, 1, 151, 5, 2, 152, 2, 14, 
/* out0467_had-eta7-phi23*/	6, 4, 0, 6, 4, 1, 8, 5, 1, 11, 5, 2, 12, 151, 4, 4, 151, 5, 14, 
/* out0468_had-eta8-phi23*/	5, 4, 0, 6, 4, 1, 7, 4, 2, 6, 151, 3, 4, 151, 4, 12, 
/* out0469_had-eta9-phi23*/	6, 3, 0, 8, 3, 1, 2, 4, 1, 1, 4, 2, 5, 150, 3, 3, 151, 3, 12, 
/* out0470_had-eta10-phi23*/	5, 3, 0, 2, 3, 1, 13, 3, 2, 5, 150, 2, 3, 150, 3, 13, 
/* out0471_had-eta11-phi23*/	5, 2, 0, 5, 2, 1, 8, 3, 1, 1, 3, 2, 4, 150, 2, 13, 
/* out0472_had-eta12-phi23*/	3, 2, 0, 2, 2, 1, 6, 2, 2, 1, 
/* out0473_had-eta13-phi23*/	4, 1, 0, 1, 1, 1, 5, 2, 1, 2, 2, 2, 5, 
/* out0474_had-eta14-phi23*/	2, 1, 0, 4, 1, 1, 3, 
/* out0475_had-eta15-phi23*/	2, 1, 1, 5, 1, 2, 1, 
/* out0476_had-eta16-phi23*/	2, 1, 1, 2, 1, 2, 3, 
/* out0477_had-eta17-phi23*/	3, 0, 0, 2, 0, 1, 2, 1, 1, 1, 
/* out0478_had-eta18-phi23*/	1, 0, 1, 6, 
/* out0479_had-eta19-phi23*/	1, 0, 1, 1, 
};