parameter integer matrixH [0:9380] = {
/* num inputs = 286(in0-in285) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 13 */
//* total number of input in adders 2966 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	1,161,0,15,
/* out0002_em-eta2-phi0*/	4,159,1,10,159,2,3,161,0,1,161,1,14,
/* out0003_em-eta3-phi0*/	7,158,0,2,158,1,15,158,2,10,159,0,5,159,1,6,160,0,15,161,1,2,
/* out0004_em-eta4-phi0*/	8,140,1,7,157,0,8,157,1,16,157,2,14,158,0,13,158,1,1,160,0,1,160,1,16,
/* out0005_em-eta5-phi0*/	10,139,1,12,139,2,6,140,0,2,140,1,1,157,0,8,157,2,2,87,0,7,87,1,15,87,2,6,94,2,3,
/* out0006_em-eta6-phi0*/	11,103,0,1,103,1,1,138,1,1,138,2,7,139,0,12,139,1,4,86,0,10,86,1,13,87,0,9,87,2,9,93,0,1,
/* out0007_em-eta7-phi0*/	11,102,1,1,102,2,1,103,0,2,138,0,8,138,1,15,138,2,9,85,0,7,85,1,3,86,0,6,86,1,1,86,2,13,
/* out0008_em-eta8-phi0*/	7,102,0,1,102,1,14,102,2,1,138,0,8,85,0,7,85,1,9,85,2,4,
/* out0009_em-eta9-phi0*/	8,101,1,1,101,2,6,102,0,7,102,1,1,84,0,1,84,1,6,85,0,2,85,2,7,
/* out0010_em-eta10-phi0*/	6,101,0,4,101,1,15,101,2,9,84,0,13,84,1,4,84,2,3,
/* out0011_em-eta11-phi0*/	8,34,1,2,34,4,3,35,1,14,101,0,6,83,0,1,83,1,4,84,0,2,84,2,5,
/* out0012_em-eta12-phi0*/	9,34,0,7,34,1,14,34,2,7,34,3,1,35,0,2,35,1,1,83,0,6,83,1,3,83,2,1,
/* out0013_em-eta13-phi0*/	7,32,5,1,33,2,2,33,5,10,34,0,9,34,3,5,83,0,3,83,2,5,
/* out0014_em-eta14-phi0*/	9,32,5,15,33,0,1,33,2,3,33,3,1,33,4,12,33,5,6,82,0,2,82,1,4,83,0,6,
/* out0015_em-eta15-phi0*/	9,32,0,6,32,1,1,32,2,16,32,3,5,33,0,15,33,3,1,33,4,4,82,0,5,82,1,1,
/* out0016_em-eta16-phi0*/	6,32,0,9,32,1,15,32,3,4,42,4,4,82,0,3,82,2,2,
/* out0017_em-eta17-phi0*/	7,32,0,1,42,4,11,43,1,1,81,0,2,81,1,2,82,0,6,82,2,1,
/* out0018_em-eta18-phi0*/	3,42,4,1,43,1,10,81,0,5,
/* out0019_em-eta19-phi0*/	3,42,1,5,43,1,2,81,0,2,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	1,161,3,15,
/* out0022_em-eta2-phi1*/	5,142,1,13,142,2,2,159,2,11,161,2,14,161,3,1,
/* out0023_em-eta3-phi1*/	10,141,0,10,141,1,14,141,2,3,142,0,3,142,1,2,158,2,5,159,0,11,159,2,2,160,3,15,161,2,2,
/* out0024_em-eta4-phi1*/	10,105,0,1,140,0,2,140,1,8,140,2,16,141,0,6,141,2,2,158,0,1,158,2,1,160,2,16,160,3,1,
/* out0025_em-eta5-phi1*/	10,104,0,5,104,1,6,139,2,7,140,0,12,87,1,1,87,2,1,93,0,2,93,1,8,94,1,14,94,2,13,
/* out0026_em-eta6-phi1*/	8,103,1,12,104,0,6,139,0,4,139,2,3,86,1,2,93,0,13,93,1,4,93,2,10,
/* out0027_em-eta7-phi1*/	8,102,2,1,103,0,13,103,1,1,103,2,6,86,2,3,92,0,12,92,1,7,92,2,1,
/* out0028_em-eta8-phi1*/	9,102,0,1,102,2,13,115,0,2,85,1,4,85,2,3,91,0,2,91,1,3,92,0,4,92,2,4,
/* out0029_em-eta9-phi1*/	5,102,0,7,114,1,6,84,1,2,85,2,2,91,0,12,
/* out0030_em-eta10-phi1*/	9,101,0,5,101,2,1,114,0,2,114,1,8,84,1,4,84,2,5,90,0,2,91,0,1,91,2,1,
/* out0031_em-eta11-phi1*/	9,34,4,13,34,5,11,35,0,5,35,1,1,101,0,1,114,0,2,83,1,3,84,2,3,90,0,6,
/* out0032_em-eta12-phi1*/	8,34,2,8,35,0,9,35,3,1,35,4,15,35,5,1,83,1,6,83,2,3,90,0,1,
/* out0033_em-eta13-phi1*/	8,33,2,1,34,2,1,34,3,10,35,3,12,35,4,1,45,1,2,83,2,7,89,0,1,
/* out0034_em-eta14-phi1*/	6,33,2,10,33,3,4,44,1,8,45,1,1,82,1,6,89,0,1,
/* out0035_em-eta15-phi1*/	6,32,3,5,33,3,10,43,5,1,44,0,4,82,1,3,82,2,3,
/* out0036_em-eta16-phi1*/	4,32,3,2,42,5,12,43,5,1,82,2,5,
/* out0037_em-eta17-phi1*/	5,42,5,4,43,0,9,43,1,1,81,1,4,82,2,1,
/* out0038_em-eta18-phi1*/	6,42,1,1,42,2,4,43,0,5,43,1,2,81,0,2,81,1,3,
/* out0039_em-eta19-phi1*/	3,42,0,1,42,1,9,81,0,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	1,163,0,15,
/* out0042_em-eta2-phi2*/	7,107,1,2,107,2,9,142,0,5,142,1,1,142,2,14,163,0,1,163,1,14,
/* out0043_em-eta3-phi2*/	8,106,0,6,106,1,16,106,2,3,141,1,2,141,2,9,142,0,8,162,0,15,163,1,2,
/* out0044_em-eta4-phi2*/	7,105,0,11,105,1,15,105,2,7,106,0,1,141,2,2,162,0,1,162,1,16,
/* out0045_em-eta5-phi2*/	11,104,0,1,104,1,10,104,2,9,105,0,4,105,2,2,117,1,3,70,0,13,70,1,9,70,2,15,93,1,2,94,1,2,
/* out0046_em-eta6-phi2*/	12,103,1,2,103,2,2,104,0,4,104,2,7,116,1,10,69,0,12,69,1,6,70,1,1,70,2,1,92,1,1,93,1,2,93,2,6,
/* out0047_em-eta7-phi2*/	10,103,2,8,115,1,7,116,0,3,116,1,3,68,0,2,68,1,1,69,0,4,69,2,2,92,1,8,92,2,6,
/* out0048_em-eta8-phi2*/	6,115,0,10,115,1,6,115,2,2,68,0,6,91,1,8,92,2,5,
/* out0049_em-eta9-phi2*/	6,114,1,1,114,2,9,115,0,4,91,0,1,91,1,5,91,2,10,
/* out0050_em-eta10-phi2*/	6,114,0,7,114,1,1,114,2,4,90,0,1,90,1,9,91,2,4,
/* out0051_em-eta11-phi2*/	7,34,5,5,35,5,5,46,4,14,114,0,4,90,0,5,90,1,2,90,2,4,
/* out0052_em-eta12-phi2*/	10,35,2,12,35,3,1,35,5,10,46,1,1,46,4,1,47,1,9,89,0,1,89,1,3,90,0,1,90,2,3,
/* out0053_em-eta13-phi2*/	7,35,2,4,35,3,2,44,4,10,45,0,1,45,1,10,89,0,7,89,1,1,
/* out0054_em-eta14-phi2*/	6,44,1,7,44,2,7,45,0,5,45,1,3,82,1,1,89,0,5,
/* out0055_em-eta15-phi2*/	7,44,0,11,44,1,1,44,2,3,44,3,5,82,1,1,82,2,2,88,0,1,
/* out0056_em-eta16-phi2*/	6,43,2,1,43,5,13,44,0,1,44,3,1,82,2,2,88,0,3,
/* out0057_em-eta17-phi2*/	5,43,0,2,43,4,11,43,5,1,81,1,3,88,0,2,
/* out0058_em-eta18-phi2*/	4,42,2,9,43,4,2,81,0,2,81,1,3,
/* out0059_em-eta19-phi2*/	5,42,0,12,42,1,1,42,2,2,42,3,1,81,0,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	1,163,3,15,
/* out0062_em-eta2-phi3*/	6,107,1,14,107,2,6,119,1,4,119,2,2,163,2,14,163,3,1,
/* out0063_em-eta3-phi3*/	9,106,0,8,106,2,13,107,2,1,118,1,3,118,2,4,119,0,4,119,1,12,162,3,15,163,2,2,
/* out0064_em-eta4-phi3*/	10,105,1,1,105,2,7,106,0,1,117,1,1,117,2,3,118,0,9,118,1,13,118,2,3,162,2,16,162,3,1,
/* out0065_em-eta5-phi3*/	7,117,0,10,117,1,12,117,2,9,70,0,3,70,1,6,73,0,11,73,1,7,
/* out0066_em-eta6-phi3*/	11,116,0,1,116,1,3,116,2,16,117,0,4,128,1,2,69,1,10,69,2,8,72,0,3,72,1,1,73,0,5,73,2,2,
/* out0067_em-eta7-phi3*/	8,115,1,2,115,2,1,116,0,12,127,1,5,68,0,1,68,1,13,69,2,6,72,0,4,
/* out0068_em-eta8-phi3*/	7,115,1,1,115,2,11,126,1,2,127,1,3,68,0,7,68,1,1,68,2,11,
/* out0069_em-eta9-phi3*/	7,114,2,1,115,2,2,126,0,5,126,1,6,67,0,8,67,1,6,91,2,1,
/* out0070_em-eta10-phi3*/	8,46,5,4,47,5,8,114,0,1,114,2,2,126,0,6,67,0,8,67,2,1,90,1,4,
/* out0071_em-eta11-phi3*/	10,46,2,1,46,4,1,46,5,12,47,0,13,47,1,1,47,4,7,47,5,5,66,0,3,90,1,1,90,2,7,
/* out0072_em-eta12-phi3*/	8,46,0,2,46,1,14,46,2,8,47,0,3,47,1,6,66,0,2,89,1,6,90,2,2,
/* out0073_em-eta13-phi3*/	9,44,4,6,44,5,14,45,0,4,45,5,1,46,0,2,46,1,1,89,0,1,89,1,4,89,2,3,
/* out0074_em-eta14-phi3*/	5,44,2,3,45,0,6,45,4,13,45,5,1,89,2,6,
/* out0075_em-eta15-phi3*/	6,44,2,3,44,3,6,45,3,7,45,4,2,88,0,1,88,1,4,
/* out0076_em-eta16-phi3*/	5,43,2,10,44,3,4,45,3,1,88,0,4,88,1,1,
/* out0077_em-eta17-phi3*/	4,43,2,4,43,3,7,43,4,2,88,0,4,
/* out0078_em-eta18-phi3*/	7,42,2,1,42,3,6,43,3,3,43,4,1,81,0,1,81,1,1,88,0,1,
/* out0079_em-eta19-phi3*/	3,0,0,1,42,0,3,42,3,5,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	1,165,0,15,
/* out0082_em-eta2-phi4*/	5,119,2,7,131,1,3,131,2,5,165,0,1,165,1,14,
/* out0083_em-eta3-phi4*/	8,118,2,3,119,0,12,119,2,7,130,0,5,130,1,12,131,2,7,164,0,15,165,1,2,
/* out0084_em-eta4-phi4*/	7,118,0,7,118,2,6,129,1,8,129,2,7,130,0,9,164,0,1,164,1,16,
/* out0085_em-eta5-phi4*/	10,117,0,2,117,2,4,128,1,2,128,2,5,129,0,8,129,1,8,73,1,9,73,2,8,74,1,5,74,2,2,
/* out0086_em-eta6-phi4*/	8,128,0,9,128,1,12,128,2,4,72,0,2,72,1,14,72,2,1,73,2,6,74,1,4,
/* out0087_em-eta7-phi4*/	9,127,0,1,127,1,6,127,2,12,128,0,2,68,1,1,68,2,1,71,1,4,72,0,7,72,2,10,
/* out0088_em-eta8-phi4*/	7,126,1,3,127,0,12,127,1,2,67,1,1,68,2,4,71,0,12,71,1,2,
/* out0089_em-eta9-phi4*/	6,126,0,1,126,1,5,126,2,8,67,1,9,67,2,6,71,0,2,
/* out0090_em-eta10-phi4*/	7,47,2,6,47,5,1,48,0,1,126,0,4,126,2,4,66,1,4,67,2,9,
/* out0091_em-eta11-phi4*/	9,46,2,1,47,2,10,47,3,14,47,4,9,47,5,2,48,0,1,66,0,5,66,1,6,66,2,1,
/* out0092_em-eta12-phi4*/	7,7,5,3,46,0,9,46,2,6,46,3,14,66,0,6,66,2,2,89,1,1,
/* out0093_em-eta13-phi4*/	8,6,5,8,7,5,5,44,5,2,45,5,7,46,0,3,60,1,2,89,1,1,89,2,4,
/* out0094_em-eta14-phi4*/	9,6,4,2,6,5,1,45,2,12,45,3,1,45,4,1,45,5,7,60,1,2,88,1,1,89,2,3,
/* out0095_em-eta15-phi4*/	5,3,2,3,3,5,4,45,2,4,45,3,7,88,1,5,
/* out0096_em-eta16-phi4*/	4,2,5,7,3,5,8,88,1,2,88,2,2,
/* out0097_em-eta17-phi4*/	5,2,4,4,2,5,6,43,2,1,43,3,2,88,2,4,
/* out0098_em-eta18-phi4*/	6,0,1,2,1,1,1,2,4,3,42,3,3,43,3,4,88,2,2,
/* out0099_em-eta19-phi4*/	3,0,0,13,0,1,8,42,3,1,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	1,165,3,15,
/* out0102_em-eta2-phi5*/	3,131,1,7,165,2,14,165,3,1,
/* out0103_em-eta3-phi5*/	7,52,1,2,130,1,4,130,2,11,131,1,6,131,2,4,164,3,15,165,2,2,
/* out0104_em-eta4-phi5*/	7,52,0,11,52,1,10,129,2,8,130,0,2,130,2,5,164,2,16,164,3,1,
/* out0105_em-eta5-phi5*/	10,51,0,13,51,1,4,51,2,1,52,0,1,128,2,2,129,0,8,129,2,1,74,0,6,74,1,2,74,2,14,
/* out0106_em-eta6-phi5*/	12,50,0,5,50,1,4,51,0,3,51,2,3,128,0,5,128,2,5,72,1,1,72,2,2,74,0,10,74,1,5,77,0,3,77,1,8,
/* out0107_em-eta7-phi5*/	6,50,0,11,50,2,4,127,2,4,71,1,6,72,2,3,77,0,13,
/* out0108_em-eta8-phi5*/	6,49,0,10,49,1,4,127,0,3,71,0,1,71,1,4,71,2,13,
/* out0109_em-eta9-phi5*/	8,48,1,1,49,0,6,49,2,4,126,2,3,71,0,1,71,2,3,75,1,4,75,2,8,
/* out0110_em-eta10-phi5*/	5,48,0,8,48,1,3,126,2,1,66,1,2,75,1,11,
/* out0111_em-eta11-phi5*/	5,47,3,2,48,0,6,48,2,3,66,1,4,66,2,6,
/* out0112_em-eta12-phi5*/	7,7,2,16,7,3,4,7,4,4,7,5,5,46,3,2,60,2,2,66,2,7,
/* out0113_em-eta13-phi5*/	6,6,5,6,7,0,11,7,4,7,7,5,3,60,1,3,60,2,5,
/* out0114_em-eta14-phi5*/	6,3,2,3,6,4,14,6,5,1,7,0,1,7,1,4,60,1,7,
/* out0115_em-eta15-phi5*/	7,3,2,10,3,3,4,3,4,3,3,5,3,60,1,2,88,1,3,88,2,1,
/* out0116_em-eta16-phi5*/	5,2,5,1,3,0,6,3,4,9,3,5,1,88,2,4,
/* out0117_em-eta17-phi5*/	5,2,4,3,2,5,2,3,0,6,3,1,2,88,2,3,
/* out0118_em-eta18-phi5*/	3,1,1,7,2,4,6,3,1,1,
/* out0119_em-eta19-phi5*/	6,0,0,2,0,1,6,0,2,12,0,3,1,1,0,4,1,1,4,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	1,167,0,15,
/* out0122_em-eta2-phi6*/	3,63,2,7,167,0,1,167,1,14,
/* out0123_em-eta3-phi6*/	7,52,1,1,62,0,11,62,1,4,63,1,4,63,2,6,166,0,15,167,1,2,
/* out0124_em-eta4-phi6*/	8,52,0,3,52,1,3,52,2,16,61,1,8,62,0,5,62,2,2,166,0,1,166,1,16,
/* out0125_em-eta5-phi6*/	10,51,1,12,51,2,6,52,0,1,60,0,1,60,1,1,61,0,8,61,1,1,79,0,6,79,1,14,79,2,2,
/* out0126_em-eta6-phi6*/	9,50,1,9,51,2,6,60,0,10,77,1,8,77,2,3,78,1,2,78,2,1,79,0,10,79,2,5,
/* out0127_em-eta7-phi6*/	6,50,1,3,50,2,12,59,1,4,76,2,6,77,2,13,78,1,3,
/* out0128_em-eta8-phi6*/	6,49,1,12,49,2,2,59,0,3,76,0,1,76,1,13,76,2,4,
/* out0129_em-eta9-phi6*/	7,48,1,1,49,2,10,58,0,3,75,0,5,75,2,8,76,0,1,76,1,3,
/* out0130_em-eta10-phi6*/	6,48,1,10,48,2,1,58,0,1,61,2,2,75,0,11,75,1,1,
/* out0131_em-eta11-phi6*/	4,19,5,2,48,2,9,61,1,6,61,2,4,
/* out0132_em-eta12-phi6*/	8,6,2,2,6,3,12,7,3,12,7,4,3,18,5,2,48,2,1,60,2,2,61,1,7,
/* out0133_em-eta13-phi6*/	8,6,0,1,6,1,5,6,2,14,6,3,2,7,0,3,7,4,2,60,0,3,60,2,6,
/* out0134_em-eta14-phi6*/	5,3,3,2,6,1,6,7,0,1,7,1,12,60,0,6,
/* out0135_em-eta15-phi6*/	7,2,2,1,2,3,6,3,3,10,3,4,2,53,1,1,53,2,3,60,0,2,
/* out0136_em-eta16-phi6*/	5,2,2,12,2,3,1,3,0,1,3,4,2,53,1,4,
/* out0137_em-eta17-phi6*/	5,2,1,3,2,2,3,3,0,3,3,1,4,53,1,3,
/* out0138_em-eta18-phi6*/	3,0,4,5,1,1,1,3,1,8,
/* out0139_em-eta19-phi6*/	6,0,2,4,0,3,15,0,4,3,0,5,1,1,0,11,1,1,3,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	1,167,3,15,
/* out0142_em-eta2-phi7*/	5,63,1,5,63,2,3,75,1,7,167,2,14,167,3,1,
/* out0143_em-eta3-phi7*/	8,62,1,12,62,2,5,63,1,7,74,1,3,75,0,12,75,1,7,166,3,15,167,2,2,
/* out0144_em-eta4-phi7*/	7,61,1,7,61,2,8,62,2,9,74,0,7,74,1,6,166,2,16,166,3,1,
/* out0145_em-eta5-phi7*/	8,60,1,8,61,0,8,61,2,8,73,0,6,79,1,2,79,2,5,80,1,8,80,2,9,
/* out0146_em-eta6-phi7*/	8,60,0,5,60,1,7,60,2,13,78,0,2,78,1,1,78,2,14,79,2,4,80,1,6,
/* out0147_em-eta7-phi7*/	9,59,0,1,59,1,12,59,2,6,60,2,2,63,1,1,63,2,1,76,2,4,78,0,7,78,1,10,
/* out0148_em-eta8-phi7*/	7,58,1,3,59,0,12,59,2,2,62,2,1,63,1,4,76,0,12,76,2,2,
/* out0149_em-eta9-phi7*/	6,58,0,8,58,1,5,58,2,1,62,1,6,62,2,9,76,0,2,
/* out0150_em-eta10-phi7*/	8,19,2,6,19,3,1,48,1,1,48,2,1,58,0,4,58,2,4,61,2,4,62,1,9,
/* out0151_em-eta11-phi7*/	9,19,0,1,19,2,10,19,3,2,19,4,9,19,5,14,48,2,1,61,0,5,61,1,1,61,2,6,
/* out0152_em-eta12-phi7*/	8,6,0,2,6,3,2,18,4,9,18,5,14,19,0,6,54,2,1,61,0,6,61,1,2,
/* out0153_em-eta13-phi7*/	8,6,0,13,6,1,2,17,2,10,18,4,3,54,1,4,54,2,1,60,0,2,60,2,1,
/* out0154_em-eta14-phi7*/	6,6,1,3,16,5,5,17,5,15,53,2,1,54,1,3,60,0,3,
/* out0155_em-eta15-phi7*/	5,2,0,2,2,3,7,16,4,3,16,5,8,53,2,5,
/* out0156_em-eta16-phi7*/	5,2,0,11,2,1,2,2,3,2,53,1,2,53,2,2,
/* out0157_em-eta17-phi7*/	5,2,0,2,2,1,9,5,2,1,5,5,2,53,1,4,
/* out0158_em-eta18-phi7*/	6,0,4,3,2,1,2,3,1,1,4,5,3,5,5,4,53,1,2,
/* out0159_em-eta19-phi7*/	4,0,4,5,0,5,9,1,0,1,4,5,1,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	1,169,0,15,
/* out0162_em-eta2-phi8*/	6,75,1,2,75,2,4,87,0,14,87,2,7,169,0,1,169,1,14,
/* out0163_em-eta3-phi8*/	9,74,1,4,74,2,3,75,0,4,75,2,12,86,0,8,86,1,13,87,0,1,168,0,15,169,1,2,
/* out0164_em-eta4-phi8*/	9,73,1,4,74,0,9,74,1,3,74,2,13,85,0,7,85,1,1,86,0,1,168,0,1,168,1,16,
/* out0165_em-eta5-phi8*/	7,73,0,9,73,1,11,73,2,11,65,0,3,65,2,7,80,0,11,80,2,7,
/* out0166_em-eta6-phi8*/	12,60,2,1,72,0,1,72,1,16,72,2,3,73,0,1,73,2,3,64,1,8,64,2,10,78,0,3,78,2,1,80,0,5,80,1,2,
/* out0167_em-eta7-phi8*/	7,59,2,5,71,1,4,72,0,12,63,0,1,63,2,13,64,1,6,78,0,4,
/* out0168_em-eta8-phi8*/	7,58,1,2,59,2,3,71,0,5,71,1,7,63,0,7,63,1,11,63,2,1,
/* out0169_em-eta9-phi8*/	7,58,1,6,58,2,5,70,1,1,71,0,2,56,1,1,62,0,8,62,2,6,
/* out0170_em-eta10-phi8*/	8,18,3,4,19,3,8,58,2,6,70,0,1,70,1,2,55,2,4,62,0,8,62,1,1,
/* out0171_em-eta11-phi8*/	10,18,0,1,18,1,1,18,2,13,18,3,12,19,0,1,19,3,5,19,4,7,55,1,7,55,2,1,61,0,3,
/* out0172_em-eta12-phi8*/	8,18,1,6,18,2,3,18,4,2,19,0,8,19,1,14,54,2,6,55,1,2,61,0,2,
/* out0173_em-eta13-phi8*/	8,17,2,6,17,3,14,17,4,4,18,4,2,19,1,1,54,0,1,54,1,3,54,2,4,
/* out0174_em-eta14-phi8*/	5,16,2,2,17,0,8,17,4,12,17,5,1,54,1,6,
/* out0175_em-eta15-phi8*/	6,16,4,7,16,5,3,17,0,6,17,1,3,53,0,1,53,2,4,
/* out0176_em-eta16-phi8*/	5,2,0,1,5,2,10,16,4,5,53,0,4,53,2,1,
/* out0177_em-eta17-phi8*/	4,5,2,4,5,4,2,5,5,7,53,0,4,
/* out0178_em-eta18-phi8*/	6,4,5,6,5,0,1,5,4,1,5,5,3,46,1,2,53,0,1,
/* out0179_em-eta19-phi8*/	3,0,5,6,4,4,3,4,5,5,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	1,169,3,15,
/* out0182_em-eta2-phi9*/	7,87,0,1,87,2,9,147,0,12,147,1,3,147,2,12,169,2,14,169,3,1,
/* out0183_em-eta3-phi9*/	9,86,0,6,86,1,3,86,2,16,145,0,2,145,1,9,147,1,4,147,2,4,168,3,15,169,2,2,
/* out0184_em-eta4-phi9*/	7,85,0,7,85,1,15,85,2,11,86,0,1,145,0,2,168,2,16,168,3,1,
/* out0185_em-eta5-phi9*/	12,73,1,1,73,2,2,84,0,9,84,1,10,84,2,1,85,0,2,85,2,4,58,2,2,59,1,2,65,0,13,65,1,15,65,2,7,
/* out0186_em-eta6-phi9*/	11,72,2,10,83,1,4,84,0,7,84,2,4,57,2,1,58,1,6,58,2,2,64,0,12,64,2,6,65,1,1,65,2,2,
/* out0187_em-eta7-phi9*/	12,71,1,3,71,2,4,72,0,3,72,2,3,83,0,4,83,1,4,57,1,6,57,2,8,63,0,2,63,2,1,64,0,4,64,1,2,
/* out0188_em-eta8-phi9*/	6,71,0,5,71,1,2,71,2,10,56,2,8,57,1,5,63,0,6,
/* out0189_em-eta9-phi9*/	6,70,1,9,70,2,1,71,0,4,56,0,1,56,1,10,56,2,5,
/* out0190_em-eta10-phi9*/	6,70,0,7,70,1,4,70,2,1,55,0,1,55,2,9,56,1,4,
/* out0191_em-eta11-phi9*/	7,18,0,14,20,3,5,21,3,5,70,0,4,55,0,5,55,1,4,55,2,2,
/* out0192_em-eta12-phi9*/	10,18,0,1,18,1,9,19,1,1,21,2,12,21,3,10,21,5,1,54,0,1,54,2,3,55,0,1,55,1,3,
/* out0193_em-eta13-phi9*/	8,16,0,3,16,2,1,16,3,14,17,3,2,21,2,4,21,5,2,54,0,7,54,2,1,
/* out0194_em-eta14-phi9*/	6,16,0,4,16,1,5,16,2,12,16,3,2,47,2,1,54,0,5,
/* out0195_em-eta15-phi9*/	7,16,1,5,16,2,1,17,0,2,17,1,12,47,1,2,47,2,1,53,0,1,
/* out0196_em-eta16-phi9*/	6,5,2,1,5,3,13,16,4,1,17,1,1,47,1,2,53,0,3,
/* out0197_em-eta17-phi9*/	5,4,2,2,5,3,1,5,4,11,46,1,2,53,0,2,
/* out0198_em-eta18-phi9*/	3,5,0,9,5,4,2,46,1,4,
/* out0199_em-eta19-phi9*/	4,4,4,12,4,5,1,5,0,2,5,1,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	1,171,0,15,
/* out0202_em-eta2-phi10*/	7,147,0,4,147,1,6,148,0,11,148,1,1,148,2,7,171,0,1,171,1,14,
/* out0203_em-eta3-phi10*/	9,145,0,4,145,1,7,145,2,15,146,2,4,147,1,3,148,1,4,148,2,9,170,0,15,171,1,2,
/* out0204_em-eta4-phi10*/	10,85,2,1,144,0,2,144,1,16,144,2,8,145,0,8,145,2,1,146,1,1,146,2,1,170,0,1,170,1,16,
/* out0205_em-eta5-phi10*/	11,84,1,6,84,2,5,143,0,4,143,1,3,144,0,12,52,1,1,52,2,1,58,0,2,58,2,8,59,0,13,59,1,14,
/* out0206_em-eta6-phi10*/	8,83,1,6,83,2,7,84,2,6,143,0,7,51,2,2,58,0,13,58,1,10,58,2,4,
/* out0207_em-eta7-phi10*/	8,82,1,1,83,0,12,83,1,2,83,2,6,51,1,3,57,0,12,57,1,1,57,2,7,
/* out0208_em-eta8-phi10*/	9,71,2,2,82,0,1,82,1,13,50,1,3,50,2,4,56,0,2,56,2,3,57,0,4,57,1,4,
/* out0209_em-eta9-phi10*/	5,70,2,6,82,0,7,49,2,2,50,1,2,56,0,12,
/* out0210_em-eta10-phi10*/	8,70,0,2,70,2,8,94,1,1,49,1,5,49,2,4,55,0,2,56,0,1,56,1,1,
/* out0211_em-eta11-phi10*/	8,20,0,13,20,1,1,20,2,5,20,3,11,70,0,2,48,2,3,49,1,3,55,0,6,
/* out0212_em-eta12-phi10*/	8,20,2,9,21,0,8,21,3,1,21,4,15,21,5,1,48,1,3,48,2,6,55,0,1,
/* out0213_em-eta13-phi10*/	8,16,0,2,20,5,10,21,0,1,21,4,1,21,5,12,29,5,1,48,1,7,54,0,1,
/* out0214_em-eta14-phi10*/	6,16,0,7,16,1,2,28,5,10,29,5,2,47,2,6,54,0,1,
/* out0215_em-eta15-phi10*/	6,5,3,1,16,1,4,28,4,11,28,5,1,47,1,3,47,2,3,
/* out0216_em-eta16-phi10*/	4,4,3,12,5,3,1,28,4,2,47,1,5,
/* out0217_em-eta17-phi10*/	6,4,1,1,4,2,9,4,3,4,46,1,1,46,2,3,47,1,1,
/* out0218_em-eta18-phi10*/	6,4,1,2,4,2,5,5,0,4,5,1,1,46,1,3,46,2,1,
/* out0219_em-eta19-phi10*/	3,4,4,1,5,1,9,46,1,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	1,171,3,15,
/* out0222_em-eta2-phi11*/	4,148,0,5,148,1,5,171,2,14,171,3,1,
/* out0223_em-eta3-phi11*/	6,146,0,15,146,1,2,146,2,11,148,1,6,170,3,15,171,2,2,
/* out0224_em-eta4-phi11*/	7,144,2,7,146,0,1,146,1,13,154,1,7,154,2,8,170,2,16,170,3,1,
/* out0225_em-eta5-phi11*/	10,143,0,1,143,1,13,143,2,4,144,0,2,144,2,1,154,1,9,52,0,7,52,1,6,52,2,15,59,0,3,
/* out0226_em-eta6-phi11*/	9,83,2,1,143,0,4,143,2,12,149,2,7,51,0,3,51,2,13,52,0,2,52,1,9,58,0,1,
/* out0227_em-eta7-phi11*/	9,82,1,1,82,2,1,83,2,2,149,1,7,149,2,9,50,2,3,51,0,5,51,1,13,51,2,1,
/* out0228_em-eta8-phi11*/	7,82,0,1,82,1,1,82,2,14,149,1,1,50,0,7,50,1,4,50,2,9,
/* out0229_em-eta9-phi11*/	7,82,0,7,82,2,1,94,2,5,49,0,1,49,2,6,50,0,2,50,1,7,
/* out0230_em-eta10-phi11*/	5,94,1,10,94,2,2,49,0,6,49,1,3,49,2,4,
/* out0231_em-eta11-phi11*/	8,20,0,3,20,1,14,21,1,2,94,1,5,48,0,1,48,2,4,49,0,1,49,1,5,
/* out0232_em-eta12-phi11*/	9,20,1,1,20,2,2,20,4,7,20,5,1,21,0,7,21,1,14,48,0,5,48,1,1,48,2,3,
/* out0233_em-eta13-phi11*/	6,20,4,9,20,5,5,29,2,7,29,5,4,48,0,3,48,1,5,
/* out0234_em-eta14-phi11*/	6,28,5,3,29,0,4,29,4,7,29,5,9,47,0,2,47,2,4,
/* out0235_em-eta15-phi11*/	6,28,4,2,28,5,2,29,0,11,29,1,4,47,0,4,47,2,1,
/* out0236_em-eta16-phi11*/	5,4,0,4,28,4,1,29,1,11,47,0,2,47,1,2,
/* out0237_em-eta17-phi11*/	4,4,0,11,4,1,1,46,2,4,47,1,1,
/* out0238_em-eta18-phi11*/	4,4,0,1,4,1,10,46,1,1,46,2,4,
/* out0239_em-eta19-phi11*/	3,4,1,2,5,1,5,46,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	1,173,0,15,
/* out0242_em-eta2-phi12*/	4,156,0,6,156,2,5,173,0,1,173,1,14,
/* out0243_em-eta3-phi12*/	6,155,0,4,155,1,7,155,2,15,156,2,8,172,0,15,173,1,2,
/* out0244_em-eta4-phi12*/	8,151,1,5,151,2,2,154,0,7,154,2,8,155,0,6,155,1,9,172,0,1,172,1,16,
/* out0245_em-eta5-phi12*/	10,150,0,1,150,1,4,150,2,13,151,1,3,154,0,9,44,0,1,44,1,5,45,0,14,45,2,8,52,0,6,
/* out0246_em-eta6-phi12*/	10,96,1,1,96,2,1,149,0,7,150,0,4,150,1,12,44,0,15,44,1,3,44,2,6,51,0,3,52,0,1,
/* out0247_em-eta7-phi12*/	8,95,2,1,96,1,2,149,0,9,149,1,7,43,0,11,43,1,5,44,2,1,51,0,5,
/* out0248_em-eta8-phi12*/	8,95,1,8,95,2,8,149,1,1,42,0,1,42,1,2,43,0,5,43,2,4,50,0,6,
/* out0249_em-eta9-phi12*/	6,94,2,6,95,1,8,42,0,12,42,1,1,49,0,1,50,0,1,
/* out0250_em-eta10-phi12*/	7,94,0,9,94,2,3,41,0,2,41,1,1,42,0,2,42,2,2,49,0,6,
/* out0251_em-eta11-phi12*/	5,31,2,9,31,3,9,94,0,5,41,0,9,49,0,1,
/* out0252_em-eta12-phi12*/	9,30,5,1,31,0,1,31,2,7,31,3,1,31,4,8,31,5,14,41,0,3,41,2,1,48,0,5,
/* out0253_em-eta13-phi12*/	7,29,2,9,29,3,4,30,4,1,30,5,12,31,5,2,40,0,5,48,0,2,
/* out0254_em-eta14-phi12*/	6,28,2,4,28,3,2,29,3,8,29,4,9,40,0,5,47,0,2,
/* out0255_em-eta15-phi12*/	7,28,0,1,28,1,5,28,2,12,28,3,1,29,0,1,40,0,1,47,0,4,
/* out0256_em-eta16-phi12*/	5,28,1,11,29,1,1,37,5,3,39,0,3,47,0,2,
/* out0257_em-eta17-phi12*/	4,36,5,9,37,5,4,39,0,3,46,2,1,
/* out0258_em-eta18-phi12*/	4,36,4,5,36,5,5,39,0,1,46,2,3,
/* out0259_em-eta19-phi12*/	2,36,4,7,46,1,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	1,173,3,15,
/* out0262_em-eta2-phi13*/	6,153,0,13,153,1,2,156,0,10,156,1,7,173,2,14,173,3,1,
/* out0263_em-eta3-phi13*/	11,152,0,3,152,1,10,152,2,14,153,0,2,153,2,3,155,0,4,155,2,1,156,1,9,156,2,3,172,3,15,173,2,2,
/* out0264_em-eta4-phi13*/	9,98,1,1,151,0,9,151,1,3,151,2,14,152,0,2,152,1,6,155,0,2,172,2,16,172,3,1,
/* out0265_em-eta5-phi13*/	11,97,2,11,150,0,4,150,2,3,151,0,7,151,1,5,38,0,14,38,1,7,38,2,2,44,1,3,45,0,2,45,2,8,
/* out0266_em-eta6-phi13*/	10,96,2,12,97,1,3,97,2,2,150,0,7,37,0,7,37,1,2,38,0,2,38,2,2,44,1,5,44,2,9,
/* out0267_em-eta7-phi13*/	8,95,2,1,96,0,6,96,1,13,96,2,1,36,0,1,37,0,7,43,1,11,43,2,4,
/* out0268_em-eta8-phi13*/	6,95,0,9,95,2,6,109,1,2,36,0,7,42,1,5,43,2,8,
/* out0269_em-eta9-phi13*/	5,95,0,7,108,2,6,42,0,1,42,1,8,42,2,8,
/* out0270_em-eta10-phi13*/	6,94,0,2,108,1,2,108,2,8,35,0,1,41,1,7,42,2,5,
/* out0271_em-eta11-phi13*/	9,30,0,4,30,2,4,30,3,16,31,3,6,31,4,2,108,1,2,41,0,2,41,1,5,41,2,4,
/* out0272_em-eta12-phi13*/	7,30,1,1,30,2,12,31,0,13,31,1,1,31,4,6,40,1,3,41,2,6,
/* out0273_em-eta13-phi13*/	8,29,3,1,30,4,14,30,5,3,31,0,2,31,1,4,39,5,2,40,0,2,40,1,5,
/* out0274_em-eta14-phi13*/	6,28,3,11,29,3,3,38,5,8,39,5,1,40,0,3,40,2,4,
/* out0275_em-eta15-phi13*/	6,28,0,12,28,3,2,37,2,1,38,4,4,39,1,2,40,2,3,
/* out0276_em-eta16-phi13*/	5,28,0,3,37,2,9,37,5,5,39,0,3,39,1,2,
/* out0277_em-eta17-phi13*/	5,36,5,1,37,0,3,37,4,7,37,5,4,39,0,4,
/* out0278_em-eta18-phi13*/	6,36,4,1,36,5,1,37,0,9,37,1,5,39,0,2,39,2,1,
/* out0279_em-eta19-phi13*/	3,36,4,3,37,1,7,39,2,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	1,175,0,15,
/* out0282_em-eta2-phi14*/	7,100,0,2,100,1,9,153,0,1,153,1,14,153,2,5,175,0,1,175,1,14,
/* out0283_em-eta3-phi14*/	7,99,1,14,99,2,11,152,0,9,152,2,2,153,2,8,174,0,15,175,1,2,
/* out0284_em-eta4-phi14*/	7,98,0,7,98,1,11,98,2,15,99,1,1,152,0,2,174,0,1,174,1,16,
/* out0285_em-eta5-phi14*/	10,97,0,16,97,1,2,97,2,3,98,0,2,98,1,4,111,2,3,32,0,6,32,1,2,38,1,9,38,2,9,
/* out0286_em-eta6-phi14*/	9,96,0,2,96,2,2,97,1,11,110,2,10,32,0,7,37,0,1,37,1,14,37,2,4,38,2,3,
/* out0287_em-eta7-phi14*/	8,96,0,8,109,2,7,110,1,3,110,2,3,31,0,3,36,1,8,37,0,1,37,2,12,
/* out0288_em-eta8-phi14*/	6,109,0,2,109,1,9,109,2,6,36,0,7,36,1,5,36,2,7,
/* out0289_em-eta9-phi14*/	8,108,0,9,108,2,1,109,1,5,35,0,4,35,1,6,36,0,1,36,2,3,42,2,1,
/* out0290_em-eta10-phi14*/	6,108,0,4,108,1,7,108,2,1,35,0,10,35,2,2,41,1,1,
/* out0291_em-eta11-phi14*/	9,30,0,10,41,2,14,108,1,4,34,0,3,34,1,1,35,0,1,35,2,1,41,1,2,41,2,3,
/* out0292_em-eta12-phi14*/	9,30,0,2,30,1,15,31,1,5,40,5,1,41,2,1,41,5,9,34,0,6,40,1,2,41,2,2,
/* out0293_em-eta13-phi14*/	8,30,4,1,31,1,6,39,2,10,39,4,1,39,5,10,34,0,1,40,1,6,40,2,1,
/* out0294_em-eta14-phi14*/	5,38,5,7,39,0,7,39,4,5,39,5,3,40,2,6,
/* out0295_em-eta15-phi14*/	6,38,4,11,38,5,1,39,0,3,39,1,5,39,1,4,40,2,2,
/* out0296_em-eta16-phi14*/	5,37,2,6,37,3,8,38,4,1,39,1,1,39,1,4,
/* out0297_em-eta17-phi14*/	4,36,2,4,37,3,1,37,4,9,39,2,4,
/* out0298_em-eta18-phi14*/	4,36,1,1,36,2,8,37,0,3,39,2,3,
/* out0299_em-eta19-phi14*/	3,36,1,5,37,0,1,37,1,4,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	1,175,3,15,
/* out0302_em-eta2-phi15*/	5,100,0,14,100,1,6,113,2,6,175,2,14,175,3,1,
/* out0303_em-eta3-phi15*/	9,99,0,15,99,2,5,100,1,1,112,0,4,112,2,3,113,1,12,113,2,4,174,3,15,175,2,2,
/* out0304_em-eta4-phi15*/	12,98,0,7,98,2,1,99,0,1,99,1,1,111,0,3,111,2,1,112,0,3,112,1,9,112,2,13,28,0,1,174,2,16,174,3,1,
/* out0305_em-eta5-phi15*/	10,111,0,9,111,1,10,111,2,12,26,0,1,28,0,10,28,1,1,28,2,16,32,0,1,32,1,14,32,2,3,
/* out0306_em-eta6-phi15*/	10,110,0,16,110,1,1,110,2,3,111,1,4,122,1,1,26,0,2,31,0,1,31,1,10,32,0,2,32,2,13,
/* out0307_em-eta7-phi15*/	9,109,0,1,109,2,2,110,1,12,121,1,2,121,2,3,31,0,12,31,1,3,31,2,7,36,1,1,
/* out0308_em-eta8-phi15*/	9,109,0,11,109,2,1,120,2,2,121,1,4,30,0,8,30,1,4,31,2,1,36,1,2,36,2,5,
/* out0309_em-eta9-phi15*/	8,108,0,1,109,0,2,120,1,5,120,2,6,30,0,6,35,1,9,35,2,1,36,2,1,
/* out0310_em-eta10-phi15*/	8,40,3,8,41,3,4,108,0,2,108,1,1,120,1,6,29,0,1,35,1,1,35,2,11,
/* out0311_em-eta11-phi15*/	10,40,2,7,40,3,5,41,0,1,41,2,1,41,3,12,41,4,13,41,5,1,34,0,1,34,1,10,35,2,1,
/* out0312_em-eta12-phi15*/	8,40,4,2,40,5,14,41,0,8,41,4,3,41,5,6,34,0,4,34,1,1,34,2,4,
/* out0313_em-eta13-phi15*/	10,38,3,1,39,2,6,39,3,14,39,4,4,40,4,2,40,5,1,33,0,1,33,1,2,34,0,1,34,2,3,
/* out0314_em-eta14-phi15*/	5,38,2,13,38,3,1,39,0,3,39,4,6,33,0,6,
/* out0315_em-eta15-phi15*/	6,38,1,7,38,2,2,39,0,3,39,1,6,33,0,5,39,1,1,
/* out0316_em-eta16-phi15*/	6,36,3,3,37,3,6,38,1,1,39,1,4,39,1,3,39,2,1,
/* out0317_em-eta17-phi15*/	4,36,2,2,36,3,11,37,3,1,39,2,4,
/* out0318_em-eta18-phi15*/	5,36,0,5,36,1,3,36,2,2,36,3,1,39,2,2,
/* out0319_em-eta19-phi15*/	3,8,3,5,36,0,2,36,1,7,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	1,177,0,15,
/* out0322_em-eta2-phi16*/	6,113,0,2,113,2,5,125,0,3,125,1,5,177,0,1,177,1,14,
/* out0323_em-eta3-phi16*/	9,112,0,3,113,0,14,113,1,4,113,2,1,124,1,5,124,2,12,125,1,7,176,0,15,177,1,2,
/* out0324_em-eta4-phi16*/	7,112,0,6,112,1,7,123,0,7,123,2,8,124,1,9,176,0,1,176,1,16,
/* out0325_em-eta5-phi16*/	12,111,0,4,111,1,2,122,2,8,123,1,8,123,2,8,26,0,1,26,1,12,27,0,2,27,1,13,27,2,1,28,0,5,28,1,15,
/* out0326_em-eta6-phi16*/	8,122,0,5,122,1,13,122,2,7,25,1,1,26,0,12,26,1,2,26,2,10,31,1,2,
/* out0327_em-eta7-phi16*/	9,121,0,5,121,1,1,121,2,13,122,1,2,25,0,11,25,1,3,30,1,1,31,1,1,31,2,8,
/* out0328_em-eta8-phi16*/	7,120,2,3,121,0,4,121,1,9,25,0,2,30,0,1,30,1,11,30,2,5,
/* out0329_em-eta9-phi16*/	6,120,0,8,120,1,1,120,2,5,29,1,5,30,0,1,30,2,9,
/* out0330_em-eta10-phi16*/	7,40,0,6,40,3,1,53,0,1,120,0,4,120,1,4,29,0,10,29,1,3,
/* out0331_em-eta11-phi16*/	10,40,0,10,40,1,14,40,2,9,40,3,2,41,0,1,53,0,1,29,0,5,29,2,1,34,1,4,34,2,1,
/* out0332_em-eta12-phi16*/	6,15,5,3,40,4,9,41,0,6,41,1,14,14,1,2,34,2,7,
/* out0333_em-eta13-phi16*/	8,14,5,8,15,5,5,38,3,7,39,3,2,40,4,3,14,1,1,33,1,6,34,2,1,
/* out0334_em-eta14-phi16*/	9,14,4,2,14,5,1,38,0,12,38,1,1,38,2,1,38,3,7,33,0,1,33,1,4,33,2,1,
/* out0335_em-eta15-phi16*/	6,13,2,2,13,3,6,38,0,4,38,1,7,33,0,2,33,2,4,
/* out0336_em-eta16-phi16*/	6,13,2,12,13,3,2,13,5,1,0,1,2,33,0,1,33,2,1,
/* out0337_em-eta17-phi16*/	5,13,2,2,13,5,8,36,0,2,36,3,1,0,1,3,
/* out0338_em-eta18-phi16*/	5,8,0,3,13,5,2,36,0,6,0,0,2,0,1,2,
/* out0339_em-eta19-phi16*/	3,8,0,5,8,3,9,36,0,1,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	1,177,3,15,
/* out0342_em-eta2-phi17*/	3,125,0,7,177,2,14,177,3,1,
/* out0343_em-eta3-phi17*/	7,57,1,1,124,0,11,124,2,4,125,0,6,125,1,4,176,3,15,177,2,2,
/* out0344_em-eta4-phi17*/	8,57,0,16,57,1,2,57,2,3,123,0,8,124,0,5,124,1,2,176,2,16,176,3,1,
/* out0345_em-eta5-phi17*/	13,56,0,13,56,1,4,56,2,1,57,2,1,122,0,1,122,2,1,123,0,1,123,1,8,23,1,5,26,1,2,27,0,14,27,1,3,27,2,15,
/* out0346_em-eta6-phi17*/	9,55,0,5,55,1,4,56,0,3,56,2,3,122,0,10,23,0,15,23,1,2,25,1,4,26,2,6,
/* out0347_em-eta7-phi17*/	6,55,0,11,55,2,4,121,0,4,25,0,2,25,1,8,25,2,13,
/* out0348_em-eta8-phi17*/	8,54,0,2,54,1,12,121,0,3,19,1,5,19,2,8,25,0,1,25,2,3,30,2,1,
/* out0349_em-eta9-phi17*/	6,53,1,1,54,0,10,120,0,3,19,1,11,29,1,5,30,2,1,
/* out0350_em-eta10-phi17*/	5,53,0,8,53,1,3,120,0,1,29,1,3,29,2,10,
/* out0351_em-eta11-phi17*/	5,40,1,2,53,0,6,53,2,3,14,2,6,29,2,5,
/* out0352_em-eta12-phi17*/	7,15,2,16,15,3,4,15,4,4,15,5,5,41,1,2,14,1,8,14,2,2,
/* out0353_em-eta13-phi17*/	6,14,5,6,15,0,11,15,4,7,15,5,3,14,1,5,33,1,2,
/* out0354_em-eta14-phi17*/	7,12,3,2,14,4,14,14,5,1,15,0,1,15,1,4,33,1,2,33,2,5,
/* out0355_em-eta15-phi17*/	5,12,2,2,12,3,9,13,3,7,13,4,1,33,2,5,
/* out0356_em-eta16-phi17*/	6,12,2,2,13,0,1,13,3,1,13,4,12,13,5,1,0,1,4,
/* out0357_em-eta17-phi17*/	5,12,5,4,13,0,3,13,4,3,13,5,4,0,1,3,
/* out0358_em-eta18-phi17*/	4,8,0,5,8,1,1,12,5,7,0,0,4,
/* out0359_em-eta19-phi17*/	6,8,0,3,8,1,3,8,2,11,8,3,2,8,5,15,9,0,2,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	1,179,0,15,
/* out0362_em-eta2-phi18*/	3,69,0,7,179,0,1,179,1,14,
/* out0363_em-eta3-phi18*/	7,57,1,2,68,0,3,68,1,12,69,0,6,69,2,4,178,0,15,179,1,2,
/* out0364_em-eta4-phi18*/	7,57,1,11,57,2,11,67,0,6,67,1,2,68,0,7,178,0,1,178,1,16,
/* out0365_em-eta5-phi18*/	12,56,1,12,56,2,6,57,2,1,66,0,1,66,1,1,67,0,8,67,2,1,21,2,2,23,1,6,24,0,15,24,1,9,24,2,16,
/* out0366_em-eta6-phi18*/	8,55,1,9,56,2,6,66,0,10,20,2,4,21,1,6,23,0,1,23,1,3,23,2,16,
/* out0367_em-eta7-phi18*/	6,55,1,3,55,2,12,65,0,4,20,0,2,20,1,13,20,2,8,
/* out0368_em-eta8-phi18*/	8,54,1,4,54,2,10,65,0,3,16,1,1,19,0,5,19,2,8,20,0,1,20,1,3,
/* out0369_em-eta9-phi18*/	8,53,1,1,54,0,4,54,2,6,64,0,1,64,1,2,15,2,5,16,1,1,19,0,11,
/* out0370_em-eta10-phi18*/	4,53,1,10,53,2,1,15,1,10,15,2,3,
/* out0371_em-eta11-phi18*/	4,27,5,2,53,2,9,14,2,6,15,1,5,
/* out0372_em-eta12-phi18*/	8,14,2,2,14,3,12,15,3,12,15,4,3,26,5,2,53,2,1,14,0,7,14,2,2,
/* out0373_em-eta13-phi18*/	8,14,0,1,14,1,5,14,2,14,14,3,2,15,0,3,15,4,2,1,2,2,14,0,5,
/* out0374_em-eta14-phi18*/	6,12,0,3,14,1,6,15,0,1,15,1,12,1,1,5,1,2,2,
/* out0375_em-eta15-phi18*/	6,12,0,9,12,1,2,12,2,3,12,3,5,0,2,1,1,1,5,
/* out0376_em-eta16-phi18*/	5,12,1,1,12,2,9,13,0,6,0,1,1,0,2,4,
/* out0377_em-eta17-phi18*/	7,12,4,3,12,5,3,13,0,6,13,1,2,0,0,2,0,1,1,0,2,3,
/* out0378_em-eta18-phi18*/	4,8,1,7,12,4,6,12,5,2,0,0,5,
/* out0379_em-eta19-phi18*/	6,8,1,4,8,2,5,8,4,2,8,5,1,9,0,14,9,1,5,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	1,179,3,15,
/* out0382_em-eta2-phi19*/	6,69,0,3,69,2,5,81,0,2,81,1,5,179,2,14,179,3,1,
/* out0383_em-eta3-phi19*/	10,68,0,1,68,1,4,68,2,12,69,2,7,80,1,3,81,0,14,81,1,1,81,2,4,178,3,15,179,2,2,
/* out0384_em-eta4-phi19*/	8,67,0,1,67,1,14,68,0,5,68,2,4,80,0,7,80,1,6,178,2,16,178,3,1,
/* out0385_em-eta5-phi19*/	11,66,1,8,67,0,1,67,2,15,79,0,6,21,0,1,21,2,12,22,0,8,22,1,16,22,2,6,24,0,1,24,1,7,
/* out0386_em-eta6-phi19*/	8,66,0,5,66,1,7,66,2,13,17,2,2,20,2,1,21,0,12,21,1,10,21,2,2,
/* out0387_em-eta7-phi19*/	9,65,0,5,65,1,13,65,2,1,66,2,2,16,2,1,17,1,8,17,2,1,20,0,11,20,2,3,
/* out0388_em-eta8-phi19*/	7,64,1,3,65,0,4,65,2,9,16,0,1,16,1,5,16,2,11,20,0,2,
/* out0389_em-eta9-phi19*/	6,64,0,3,64,1,10,64,2,1,15,2,5,16,0,1,16,1,9,
/* out0390_em-eta10-phi19*/	7,27,2,6,27,3,1,53,1,1,53,2,1,64,0,9,15,0,10,15,2,3,
/* out0391_em-eta11-phi19*/	10,27,0,1,27,2,10,27,3,2,27,4,9,27,5,14,53,2,1,2,1,1,2,2,4,15,0,5,15,1,1,
/* out0392_em-eta12-phi19*/	7,14,0,2,14,3,2,26,4,9,26,5,14,27,0,6,2,1,7,14,0,3,
/* out0393_em-eta13-phi19*/	7,14,0,13,14,1,2,23,2,10,26,4,3,1,2,6,2,1,1,14,0,1,
/* out0394_em-eta14-phi19*/	6,14,1,3,22,5,5,23,5,15,1,0,1,1,1,1,1,2,4,
/* out0395_em-eta15-phi19*/	6,12,0,4,12,1,5,22,4,3,22,5,8,1,0,2,1,1,4,
/* out0396_em-eta16-phi19*/	5,12,1,8,13,1,7,0,2,3,1,0,1,1,1,1,
/* out0397_em-eta17-phi19*/	5,11,2,2,11,3,1,12,4,4,13,1,6,0,2,4,
/* out0398_em-eta18-phi19*/	6,8,1,1,9,1,3,11,2,6,12,4,3,0,0,3,0,2,1,
/* out0399_em-eta19-phi19*/	3,8,4,12,9,1,8,11,2,1,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	1,181,0,15,
/* out0402_em-eta2-phi20*/	5,81,1,6,93,0,14,93,2,6,181,0,1,181,1,14,
/* out0403_em-eta3-phi20*/	9,80,1,4,80,2,3,81,1,4,81,2,12,92,0,15,92,1,5,93,2,1,180,0,15,181,1,2,
/* out0404_em-eta4-phi20*/	11,79,1,4,80,0,9,80,1,3,80,2,13,91,0,2,91,1,5,92,0,1,92,2,1,22,2,1,180,0,1,180,1,16,
/* out0405_em-eta5-phi20*/	9,79,0,9,79,1,11,79,2,11,18,0,1,18,1,3,18,2,14,21,0,1,22,0,8,22,2,9,
/* out0406_em-eta6-phi20*/	11,66,2,1,78,0,9,78,1,10,78,2,1,79,0,1,79,2,3,17,0,1,17,2,10,18,0,2,18,1,13,21,0,2,
/* out0407_em-eta7-phi20*/	10,65,1,3,65,2,2,77,0,1,77,1,2,78,0,7,78,2,5,4,2,1,17,0,12,17,1,7,17,2,3,
/* out0408_em-eta8-phi20*/	10,64,1,1,64,2,1,65,2,4,77,0,11,77,1,1,4,1,5,4,2,2,16,0,8,16,2,4,17,1,1,
/* out0409_em-eta9-phi20*/	7,64,2,11,76,0,1,77,0,2,3,1,1,3,2,9,4,1,1,16,0,6,
/* out0410_em-eta10-phi20*/	8,26,3,4,27,3,8,64,0,3,64,2,3,76,0,3,3,1,11,3,2,1,15,0,1,
/* out0411_em-eta11-phi20*/	10,26,0,1,26,1,1,26,2,13,26,3,12,27,0,1,27,3,5,27,4,7,2,0,1,2,2,10,3,1,1,
/* out0412_em-eta12-phi20*/	8,26,1,6,26,2,3,26,4,2,27,0,8,27,1,14,2,0,4,2,1,4,2,2,1,
/* out0413_em-eta13-phi20*/	9,23,2,6,23,3,14,23,4,4,26,4,2,27,1,1,1,0,1,1,2,2,2,0,1,2,1,3,
/* out0414_em-eta14-phi20*/	5,22,2,2,23,0,8,23,4,12,23,5,1,1,0,6,
/* out0415_em-eta15-phi20*/	6,22,4,7,22,5,3,23,0,6,23,1,3,1,0,5,7,2,1,
/* out0416_em-eta16-phi20*/	6,10,3,6,11,3,3,13,1,1,22,4,5,7,1,1,7,2,3,
/* out0417_em-eta17-phi20*/	4,10,3,1,11,3,11,11,4,2,7,1,4,
/* out0418_em-eta18-phi20*/	5,11,2,5,11,3,1,11,4,2,11,5,3,7,1,2,
/* out0419_em-eta19-phi20*/	3,8,4,2,11,2,2,11,5,7,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	1,181,3,15,
/* out0422_em-eta2-phi21*/	7,93,0,2,93,2,9,137,0,12,137,1,3,137,2,12,181,2,14,181,3,1,
/* out0423_em-eta3-phi21*/	8,92,1,11,92,2,14,135,0,9,135,1,2,137,1,4,137,2,4,180,3,15,181,2,2,
/* out0424_em-eta4-phi21*/	7,91,0,8,91,1,11,91,2,15,92,2,1,135,0,2,180,2,16,180,3,1,
/* out0425_em-eta5-phi21*/	10,79,1,1,79,2,2,90,0,9,90,1,10,90,2,1,91,0,6,6,1,9,6,2,9,18,0,6,18,2,2,
/* out0426_em-eta6-phi21*/	11,78,1,6,78,2,4,89,0,2,89,1,2,90,0,7,90,2,4,5,0,1,5,1,4,5,2,14,6,1,3,18,0,7,
/* out0427_em-eta7-phi21*/	7,77,1,7,78,2,6,89,0,8,4,2,8,5,0,1,5,1,12,17,0,3,
/* out0428_em-eta8-phi21*/	6,77,0,2,77,1,6,77,2,9,4,0,7,4,1,7,4,2,5,
/* out0429_em-eta9-phi21*/	8,76,0,2,76,1,8,77,2,5,3,0,4,3,2,6,4,0,1,4,1,3,10,1,1,
/* out0430_em-eta10-phi21*/	6,76,0,8,76,1,1,76,2,2,3,0,10,3,1,2,9,2,1,
/* out0431_em-eta11-phi21*/	10,25,2,10,26,0,14,76,0,2,76,2,2,2,0,3,2,2,1,3,0,1,3,1,1,9,1,3,9,2,2,
/* out0432_em-eta12-phi21*/	9,24,5,5,25,2,2,25,5,15,26,0,1,26,1,9,27,1,1,2,0,6,8,2,2,9,1,2,
/* out0433_em-eta13-phi21*/	9,22,0,3,22,2,1,22,3,15,23,3,2,24,4,1,24,5,6,2,0,1,8,1,1,8,2,6,
/* out0434_em-eta14-phi21*/	5,22,0,4,22,1,5,22,2,12,22,3,1,8,1,6,
/* out0435_em-eta15-phi21*/	6,22,1,5,22,2,1,23,0,2,23,1,12,7,2,4,8,1,2,
/* out0436_em-eta16-phi21*/	5,10,0,6,10,3,8,22,4,1,23,1,1,7,2,4,
/* out0437_em-eta17-phi21*/	4,10,2,9,10,3,1,11,4,4,7,1,4,
/* out0438_em-eta18-phi21*/	4,11,0,3,11,4,8,11,5,1,7,1,3,
/* out0439_em-eta19-phi21*/	3,10,5,4,11,0,1,11,5,5,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	1,183,0,15,
/* out0442_em-eta2-phi22*/	6,136,0,13,136,1,6,137,0,4,137,1,6,183,0,1,183,1,14,
/* out0443_em-eta3-phi22*/	10,134,1,4,134,2,1,135,0,3,135,1,14,135,2,10,136,0,3,136,2,12,137,1,3,182,0,15,183,1,2,
/* out0444_em-eta4-phi22*/	9,91,2,1,133,0,9,133,1,14,133,2,3,134,1,2,135,0,2,135,2,6,182,0,1,182,1,16,
/* out0445_em-eta5-phi22*/	12,90,1,6,90,2,5,132,0,4,132,1,3,133,0,7,133,2,5,6,0,14,6,1,2,6,2,7,12,2,3,13,0,2,13,1,8,
/* out0446_em-eta6-phi22*/	9,89,1,12,90,2,6,132,0,7,5,0,7,5,2,2,6,0,2,6,1,2,12,1,9,12,2,5,
/* out0447_em-eta7-phi22*/	8,88,1,1,89,0,6,89,1,1,89,2,13,4,0,1,5,0,7,11,1,4,11,2,11,
/* out0448_em-eta8-phi22*/	6,77,2,2,88,0,9,88,1,6,4,0,7,10,2,5,11,1,8,
/* out0449_em-eta9-phi22*/	5,76,1,6,88,0,7,10,0,1,10,1,8,10,2,8,
/* out0450_em-eta10-phi22*/	5,76,1,1,76,2,10,3,0,1,9,2,7,10,1,5,
/* out0451_em-eta11-phi22*/	9,24,2,2,24,3,6,25,2,4,25,3,16,25,4,4,76,2,2,9,0,2,9,1,4,9,2,5,
/* out0452_em-eta12-phi22*/	7,24,2,6,24,5,1,25,0,13,25,4,12,25,5,1,8,2,3,9,1,6,
/* out0453_em-eta13-phi22*/	7,22,0,2,24,4,14,24,5,4,25,0,2,25,1,3,8,0,2,8,2,5,
/* out0454_em-eta14-phi22*/	4,22,0,7,22,1,2,8,0,3,8,1,4,
/* out0455_em-eta15-phi22*/	4,10,0,1,22,1,4,7,2,2,8,1,3,
/* out0456_em-eta16-phi22*/	4,10,0,9,10,1,5,7,0,3,7,2,2,
/* out0457_em-eta17-phi22*/	5,10,1,4,10,2,7,11,0,3,11,1,1,7,0,4,
/* out0458_em-eta18-phi22*/	6,10,4,1,10,5,5,11,0,9,11,1,1,7,0,2,7,1,1,
/* out0459_em-eta19-phi22*/	3,10,4,3,10,5,7,7,1,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	1,183,3,15,
/* out0462_em-eta2-phi23*/	3,136,1,7,183,2,14,183,3,1,
/* out0463_em-eta3-phi23*/	7,134,0,7,134,1,4,134,2,15,136,1,3,136,2,4,182,3,15,183,2,2,
/* out0464_em-eta4-phi23*/	6,133,1,2,133,2,5,134,0,9,134,1,6,182,2,16,182,3,1,
/* out0465_em-eta5-phi23*/	8,132,0,1,132,1,13,132,2,4,133,2,3,12,0,1,12,2,5,13,0,14,13,1,8,
/* out0466_em-eta6-phi23*/	7,89,1,1,89,2,1,132,0,4,132,2,12,12,0,15,12,1,6,12,2,3,
/* out0467_em-eta7-phi23*/	5,88,1,1,89,2,2,11,0,11,11,2,5,12,1,1,
/* out0468_em-eta8-phi23*/	6,88,1,8,88,2,8,10,0,1,10,2,2,11,0,5,11,1,4,
/* out0469_em-eta9-phi23*/	3,88,2,8,10,0,12,10,2,1,
/* out0470_em-eta10-phi23*/	4,9,0,2,9,2,1,10,0,2,10,1,2,
/* out0471_em-eta11-phi23*/	3,24,0,9,24,3,9,9,0,9,
/* out0472_em-eta12-phi23*/	8,24,0,7,24,1,14,24,2,8,24,3,1,25,0,1,25,1,1,9,0,3,9,1,1,
/* out0473_em-eta13-phi23*/	4,24,1,2,24,4,1,25,1,12,8,0,5,
/* out0474_em-eta14-phi23*/	1,8,0,5,
/* out0475_em-eta15-phi23*/	1,8,0,1,
/* out0476_em-eta16-phi23*/	2,10,1,3,7,0,3,
/* out0477_em-eta17-phi23*/	3,10,1,4,11,1,9,7,0,3,
/* out0478_em-eta18-phi23*/	3,10,4,5,11,1,5,7,0,1,
/* out0479_em-eta19-phi23*/	1,10,4,7
};