parameter integer matrixH [0:8348] = {
/* num inputs = 140(in0-in139) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 15 */
//* total number of input in adders 2622 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	3,79,0,7,79,1,1,89,2,2,
/* out0005_em-eta5-phi0*/	7,75,1,1,85,1,8,85,2,15,79,0,9,79,1,14,79,2,9,89,2,1,
/* out0006_em-eta6-phi0*/	9,75,0,14,75,1,7,75,2,3,68,0,16,68,1,9,68,2,2,79,2,7,80,0,1,80,2,1,
/* out0007_em-eta7-phi0*/	8,65,0,6,65,1,6,75,0,2,75,2,4,57,0,11,57,1,1,68,1,3,68,2,14,
/* out0008_em-eta8-phi0*/	6,54,1,1,65,0,10,65,2,4,57,0,5,57,1,6,57,2,8,
/* out0009_em-eta9-phi0*/	5,54,0,11,54,1,2,46,0,10,46,1,1,57,2,5,
/* out0010_em-eta10-phi0*/	7,43,0,1,43,1,1,54,0,5,54,2,2,46,0,3,46,1,3,46,2,8,
/* out0011_em-eta11-phi0*/	4,43,0,8,131,2,10,35,0,7,46,2,4,
/* out0012_em-eta12-phi0*/	9,43,0,5,43,2,1,124,0,3,124,1,2,131,1,2,131,2,2,35,0,5,35,1,1,35,2,4,
/* out0013_em-eta13-phi0*/	4,32,0,3,124,0,9,24,0,1,35,2,7,
/* out0014_em-eta14-phi0*/	5,32,0,6,117,0,1,124,0,2,124,2,1,24,0,7,
/* out0015_em-eta15-phi0*/	4,32,0,2,117,0,5,24,0,2,24,2,4,
/* out0016_em-eta16-phi0*/	3,22,0,2,117,0,4,24,2,5,
/* out0017_em-eta17-phi0*/	5,22,0,3,111,2,1,117,0,1,14,2,5,24,2,1,
/* out0018_em-eta18-phi0*/	4,22,0,1,111,2,3,14,0,1,14,2,3,
/* out0019_em-eta19-phi0*/	2,111,0,1,14,0,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	2,89,1,3,89,2,8,
/* out0025_em-eta5-phi1*/	10,85,1,8,85,2,1,86,0,11,86,1,7,86,2,1,79,1,1,80,0,14,80,1,4,89,1,11,89,2,5,
/* out0026_em-eta6-phi1*/	11,75,1,8,75,2,6,76,0,4,76,1,2,86,0,5,86,2,4,68,1,3,69,0,5,80,0,1,80,1,2,80,2,15,
/* out0027_em-eta7-phi1*/	8,65,1,10,75,2,3,76,0,11,57,1,1,68,1,1,69,0,10,69,1,1,69,2,9,
/* out0028_em-eta8-phi1*/	6,54,1,2,65,2,12,66,0,6,57,1,7,58,0,8,69,2,4,
/* out0029_em-eta9-phi1*/	9,54,1,11,54,2,4,66,0,1,46,0,3,46,1,4,57,1,1,57,2,3,58,0,3,58,2,8,
/* out0030_em-eta10-phi1*/	7,43,1,4,54,2,9,55,0,1,46,1,8,46,2,3,47,0,4,58,2,1,
/* out0031_em-eta11-phi1*/	10,43,0,1,43,1,8,43,2,2,131,1,9,131,2,4,35,0,4,35,1,3,46,2,1,47,0,2,47,2,3,
/* out0032_em-eta12-phi1*/	8,32,1,1,43,0,1,43,2,8,124,1,9,131,1,4,132,0,1,35,1,9,35,2,2,
/* out0033_em-eta13-phi1*/	10,32,0,1,32,1,7,124,0,2,124,1,3,124,2,5,24,0,1,35,1,2,35,2,3,36,0,1,36,2,1,
/* out0034_em-eta14-phi1*/	7,32,0,3,32,1,1,32,2,2,117,1,4,124,2,5,24,0,4,24,1,4,
/* out0035_em-eta15-phi1*/	8,22,1,1,32,0,1,32,2,4,117,0,3,117,1,5,24,0,1,24,1,5,24,2,1,
/* out0036_em-eta16-phi1*/	7,22,0,2,22,1,3,117,0,2,117,2,4,14,2,1,24,1,1,24,2,4,
/* out0037_em-eta17-phi1*/	6,22,0,4,111,2,4,117,2,2,14,0,1,14,2,4,24,2,1,
/* out0038_em-eta18-phi1*/	6,22,0,3,22,2,1,111,0,2,111,2,4,14,0,3,14,2,1,
/* out0039_em-eta19-phi1*/	4,22,0,1,22,2,1,111,0,1,14,0,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	3,89,1,2,90,0,5,90,1,4,
/* out0045_em-eta5-phi2*/	12,86,1,9,86,2,5,87,0,2,87,1,2,94,0,14,94,1,13,94,2,12,80,1,5,81,0,3,90,0,11,90,1,5,90,2,15,
/* out0046_em-eta6-phi2*/	8,76,1,12,86,2,6,87,0,10,69,0,1,69,1,2,80,1,5,81,0,11,81,2,8,
/* out0047_em-eta7-phi2*/	9,66,1,3,76,0,1,76,1,2,76,2,16,77,0,3,69,1,13,69,2,1,70,0,5,81,2,2,
/* out0048_em-eta8-phi2*/	8,66,0,6,66,1,10,66,2,4,58,0,5,58,1,7,69,2,2,70,0,1,70,2,3,
/* out0049_em-eta9-phi2*/	7,54,2,1,55,0,2,55,1,5,66,0,3,66,2,6,58,1,7,58,2,7,
/* out0050_em-eta10-phi2*/	5,55,0,11,55,1,2,55,2,1,47,0,9,47,1,3,
/* out0051_em-eta11-phi2*/	12,43,1,3,43,2,2,44,0,1,44,1,1,55,0,2,55,2,2,131,1,1,132,0,6,132,1,7,47,0,1,47,1,1,47,2,9,
/* out0052_em-eta12-phi2*/	8,43,2,3,44,0,7,124,1,1,132,0,9,132,2,2,35,1,1,36,0,6,47,2,2,
/* out0053_em-eta13-phi2*/	9,32,1,6,44,0,2,124,1,1,124,2,4,125,0,4,125,1,1,132,2,1,36,0,4,36,2,3,
/* out0054_em-eta14-phi2*/	7,32,1,1,32,2,6,117,1,2,124,2,1,125,0,6,24,1,2,36,2,4,
/* out0055_em-eta15-phi2*/	7,22,1,2,32,2,3,33,0,1,117,1,5,117,2,2,24,1,3,25,0,2,
/* out0056_em-eta16-phi2*/	5,22,1,5,117,2,6,14,2,1,24,1,1,25,0,2,
/* out0057_em-eta17-phi2*/	8,22,1,1,22,2,2,111,0,2,111,2,3,117,2,1,14,0,3,14,2,1,25,2,1,
/* out0058_em-eta18-phi2*/	4,22,2,3,111,0,5,111,2,1,14,0,4,
/* out0059_em-eta19-phi2*/	1,22,2,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	2,90,1,1,91,0,2,
/* out0065_em-eta5-phi3*/	13,87,1,11,94,0,2,94,1,3,94,2,4,95,0,16,95,1,4,95,2,8,81,0,1,81,1,2,90,1,6,90,2,1,91,0,13,91,2,8,
/* out0066_em-eta6-phi3*/	10,77,1,5,87,0,4,87,1,3,87,2,16,88,0,3,81,0,1,81,1,14,81,2,4,82,0,5,91,2,2,
/* out0067_em-eta7-phi3*/	7,77,0,11,77,1,8,77,2,5,70,0,10,70,1,8,81,2,2,82,2,1,
/* out0068_em-eta8-phi3*/	10,66,1,3,66,2,4,67,0,5,67,1,4,77,0,2,77,2,3,58,1,1,59,0,3,70,1,2,70,2,12,
/* out0069_em-eta9-phi3*/	6,55,1,5,66,2,2,67,0,9,58,1,1,59,0,11,59,2,4,
/* out0070_em-eta10-phi3*/	6,55,1,4,55,2,9,56,0,1,47,1,6,48,0,1,59,2,5,
/* out0071_em-eta11-phi3*/	11,44,1,7,55,2,4,56,0,1,132,1,9,132,2,2,137,0,10,137,1,7,137,2,3,47,1,6,47,2,2,48,0,3,
/* out0072_em-eta12-phi3*/	9,44,0,4,44,1,3,44,2,3,125,1,1,132,2,11,133,0,1,36,0,4,36,1,4,48,2,1,
/* out0073_em-eta13-phi3*/	8,33,1,1,44,0,2,44,2,4,125,0,1,125,1,10,36,0,1,36,1,4,36,2,2,
/* out0074_em-eta14-phi3*/	7,32,2,1,33,0,5,33,1,2,125,0,4,125,2,4,25,0,1,36,2,5,
/* out0075_em-eta15-phi3*/	7,33,0,5,117,2,1,118,0,1,118,1,3,125,0,1,125,2,2,25,0,5,
/* out0076_em-eta16-phi3*/	5,22,1,3,33,0,1,118,0,6,25,0,3,25,2,2,
/* out0077_em-eta17-phi3*/	5,22,1,1,22,2,4,111,0,1,118,0,4,25,2,3,
/* out0078_em-eta18-phi3*/	4,22,2,3,111,0,4,14,0,2,25,2,1,
/* out0079_em-eta19-phi3*/	1,22,2,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	5,91,0,1,91,1,1,97,0,11,97,1,5,97,2,8,
/* out0085_em-eta5-phi4*/	13,88,1,6,95,1,12,95,2,8,96,0,13,96,1,1,96,2,2,91,1,15,91,2,5,92,0,8,92,2,2,97,0,4,97,1,8,97,2,4,
/* out0086_em-eta6-phi4*/	8,88,0,12,88,1,8,88,2,8,82,0,11,82,1,11,82,2,3,91,2,1,92,2,1,
/* out0087_em-eta7-phi4*/	9,77,1,3,77,2,7,78,0,8,78,1,4,88,0,1,88,2,2,70,1,4,71,0,7,82,2,11,
/* out0088_em-eta8-phi4*/	10,67,1,12,67,2,2,77,2,1,78,0,5,59,0,1,59,1,3,70,1,2,70,2,1,71,0,5,71,2,6,
/* out0089_em-eta9-phi4*/	6,56,1,2,67,0,2,67,2,12,59,0,1,59,1,12,59,2,2,
/* out0090_em-eta10-phi4*/	6,56,0,7,56,1,6,48,0,6,48,1,1,59,1,1,59,2,5,
/* out0091_em-eta11-phi4*/	11,44,1,3,56,0,7,56,2,1,133,0,1,133,1,6,137,0,6,137,1,9,137,2,13,48,0,6,48,1,1,48,2,4,
/* out0092_em-eta12-phi4*/	8,44,1,2,44,2,6,45,0,2,133,0,11,133,1,2,133,2,1,36,1,2,48,2,6,
/* out0093_em-eta13-phi4*/	10,33,1,3,44,2,3,45,0,1,125,1,4,125,2,2,126,0,1,133,0,3,133,2,1,36,1,5,37,0,3,
/* out0094_em-eta14-phi4*/	10,33,0,1,33,1,6,125,2,7,126,0,2,25,0,1,25,1,1,36,1,1,36,2,1,37,0,1,37,2,1,
/* out0095_em-eta15-phi4*/	6,33,0,2,33,2,3,118,1,6,125,2,1,25,0,2,25,1,4,
/* out0096_em-eta16-phi4*/	8,23,2,1,33,0,1,33,2,2,118,0,2,118,1,3,118,2,2,25,1,2,25,2,2,
/* out0097_em-eta17-phi4*/	4,23,1,3,118,0,2,118,2,3,25,2,4,
/* out0098_em-eta18-phi4*/	4,23,1,3,118,0,1,118,2,1,25,2,1,
/* out0099_em-eta19-phi4*/	0,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	6,97,0,1,97,1,2,97,2,3,98,0,5,98,1,1,98,2,3,
/* out0105_em-eta5-phi5*/	12,89,1,2,96,0,3,96,1,15,96,2,13,92,0,8,92,1,16,92,2,6,97,1,1,97,2,1,98,0,7,98,1,7,98,2,1,
/* out0106_em-eta6-phi5*/	9,88,1,2,88,2,6,89,0,14,89,1,6,96,2,1,82,1,4,83,0,15,83,2,1,92,2,7,
/* out0107_em-eta7-phi5*/	10,78,0,1,78,1,12,78,2,8,89,0,2,71,0,3,71,1,9,82,1,1,82,2,1,83,0,1,83,2,7,
/* out0108_em-eta8-phi5*/	9,67,2,1,68,0,2,68,1,7,78,0,2,78,2,8,60,0,2,71,0,1,71,1,7,71,2,9,
/* out0109_em-eta9-phi5*/	7,56,1,2,67,2,1,68,0,13,68,1,1,60,0,13,60,2,1,71,2,1,
/* out0110_em-eta10-phi5*/	6,56,1,6,56,2,7,68,0,1,48,1,5,60,0,1,60,2,7,
/* out0111_em-eta11-phi5*/	8,45,1,3,56,2,8,133,1,6,138,0,12,138,1,8,138,2,4,48,1,9,48,2,1,
/* out0112_em-eta12-phi5*/	6,45,0,5,45,1,5,133,1,2,133,2,11,37,0,4,48,2,4,
/* out0113_em-eta13-phi5*/	6,33,1,1,45,0,7,126,0,1,126,1,7,133,2,3,37,0,7,
/* out0114_em-eta14-phi5*/	7,33,1,3,33,2,3,45,0,1,126,0,8,126,1,1,37,0,1,37,2,6,
/* out0115_em-eta15-phi5*/	5,33,2,6,118,1,3,126,0,4,25,1,4,37,2,1,
/* out0116_em-eta16-phi5*/	5,23,2,4,33,2,2,118,1,1,118,2,5,25,1,4,
/* out0117_em-eta17-phi5*/	5,23,1,1,23,2,2,118,2,5,25,1,1,25,2,2,
/* out0118_em-eta18-phi5*/	1,23,1,3,
/* out0119_em-eta19-phi5*/	1,23,1,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	6,98,0,3,98,1,1,98,2,5,99,0,3,99,1,2,99,2,1,
/* out0125_em-eta5-phi6*/	12,89,1,2,97,0,16,97,1,11,97,2,13,93,0,16,93,1,8,93,2,6,98,0,1,98,1,7,98,2,7,99,0,1,99,1,1,
/* out0126_em-eta6-phi6*/	9,89,1,6,89,2,14,90,0,6,90,1,2,97,2,1,83,1,15,83,2,1,84,0,4,93,2,7,
/* out0127_em-eta7-phi6*/	10,79,0,8,79,1,12,79,2,1,89,2,2,72,0,9,72,1,3,83,1,1,83,2,7,84,0,1,84,2,1,
/* out0128_em-eta8-phi6*/	9,68,1,7,68,2,2,69,0,1,79,0,8,79,2,2,60,1,2,72,0,7,72,1,1,72,2,9,
/* out0129_em-eta9-phi6*/	7,57,1,2,68,1,1,68,2,13,69,0,1,60,1,13,60,2,1,72,2,1,
/* out0130_em-eta10-phi6*/	6,57,0,7,57,1,6,68,2,1,49,0,5,60,1,1,60,2,7,
/* out0131_em-eta11-phi6*/	8,45,1,3,57,0,8,134,1,6,138,0,4,138,1,8,138,2,12,49,0,9,49,2,1,
/* out0132_em-eta12-phi6*/	6,45,1,5,45,2,5,134,0,11,134,1,2,37,1,4,49,2,4,
/* out0133_em-eta13-phi6*/	6,34,1,1,45,2,7,126,1,7,126,2,1,134,0,3,37,1,7,
/* out0134_em-eta14-phi6*/	7,34,0,3,34,1,3,45,2,1,126,1,1,126,2,8,37,1,1,37,2,6,
/* out0135_em-eta15-phi6*/	5,34,0,6,119,1,3,126,2,4,26,0,4,37,2,1,
/* out0136_em-eta16-phi6*/	5,23,2,4,34,0,2,119,0,5,119,1,1,26,0,4,
/* out0137_em-eta17-phi6*/	5,23,0,2,23,2,3,119,0,5,26,0,1,26,2,2,
/* out0138_em-eta18-phi6*/	2,23,0,1,23,1,3,
/* out0139_em-eta19-phi6*/	1,23,1,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	5,94,0,1,94,1,1,99,0,8,99,1,5,99,2,11,
/* out0145_em-eta5-phi7*/	13,90,1,6,97,1,5,97,2,2,98,0,16,98,1,7,98,2,8,93,1,8,93,2,2,94,0,15,94,2,5,99,0,4,99,1,8,99,2,4,
/* out0146_em-eta6-phi7*/	8,90,0,8,90,1,8,90,2,12,84,0,11,84,1,11,84,2,3,93,2,1,94,2,1,
/* out0147_em-eta7-phi7*/	9,79,1,4,79,2,8,80,0,7,80,1,3,90,0,2,90,2,1,72,1,7,73,0,4,84,2,11,
/* out0148_em-eta8-phi7*/	10,69,0,2,69,1,12,79,2,5,80,0,1,61,0,3,61,1,1,72,1,5,72,2,6,73,0,2,73,2,1,
/* out0149_em-eta9-phi7*/	6,57,1,2,69,0,12,69,2,2,61,0,12,61,1,1,61,2,2,
/* out0150_em-eta10-phi7*/	6,57,1,6,57,2,7,49,0,1,49,1,6,61,0,1,61,2,5,
/* out0151_em-eta11-phi7*/	11,46,1,3,57,0,1,57,2,7,134,1,6,134,2,1,139,0,13,139,1,9,139,2,6,49,0,1,49,1,6,49,2,4,
/* out0152_em-eta12-phi7*/	8,45,2,2,46,0,6,46,1,2,134,0,1,134,1,2,134,2,11,38,0,2,49,2,6,
/* out0153_em-eta13-phi7*/	10,34,1,3,45,2,1,46,0,3,126,2,1,127,0,2,127,1,4,134,0,1,134,2,3,37,1,3,38,0,5,
/* out0154_em-eta14-phi7*/	10,34,1,6,34,2,1,126,2,2,127,0,7,26,0,1,26,1,1,37,1,1,37,2,1,38,0,1,38,2,1,
/* out0155_em-eta15-phi7*/	6,34,0,3,34,2,2,119,1,6,127,0,1,26,0,4,26,1,2,
/* out0156_em-eta16-phi7*/	8,23,2,1,34,0,2,34,2,1,119,0,2,119,1,3,119,2,2,26,0,2,26,2,2,
/* out0157_em-eta17-phi7*/	5,23,0,7,23,2,1,119,0,3,119,2,2,26,2,4,
/* out0158_em-eta18-phi7*/	5,23,0,5,23,1,1,119,0,1,119,2,1,26,2,1,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	2,94,1,2,95,1,1,
/* out0165_em-eta5-phi8*/	13,91,1,11,98,1,9,98,2,8,99,0,4,99,1,3,99,2,2,85,0,2,85,1,1,94,1,13,94,2,8,95,0,13,95,1,1,95,2,1,
/* out0166_em-eta6-phi8*/	10,80,1,5,90,2,3,91,0,16,91,1,3,91,2,4,84,1,5,85,0,14,85,1,1,85,2,4,94,2,2,
/* out0167_em-eta7-phi8*/	7,80,0,5,80,1,8,80,2,11,73,0,8,73,1,10,84,2,1,85,2,2,
/* out0168_em-eta8-phi8*/	10,69,1,4,69,2,5,70,0,4,70,1,3,80,0,3,80,2,2,61,1,3,62,0,1,73,0,2,73,2,12,
/* out0169_em-eta9-phi8*/	6,58,1,5,69,2,9,70,0,2,61,1,11,61,2,4,62,0,1,
/* out0170_em-eta10-phi8*/	6,57,2,1,58,0,9,58,1,4,49,1,1,50,0,6,61,2,5,
/* out0171_em-eta11-phi8*/	11,46,1,7,57,2,1,58,0,4,135,0,2,135,1,9,139,0,3,139,1,7,139,2,10,49,1,3,50,0,6,50,2,2,
/* out0172_em-eta12-phi8*/	9,46,0,3,46,1,3,46,2,4,127,1,1,134,2,1,135,0,11,38,0,4,38,1,4,49,2,1,
/* out0173_em-eta13-phi8*/	8,34,1,1,46,0,4,46,2,2,127,1,10,127,2,1,38,0,4,38,1,1,38,2,2,
/* out0174_em-eta14-phi8*/	7,34,1,2,34,2,5,35,0,1,127,0,4,127,2,4,26,1,1,38,2,5,
/* out0175_em-eta15-phi8*/	7,34,2,5,119,1,3,119,2,1,120,0,1,127,0,2,127,2,1,26,1,5,
/* out0176_em-eta16-phi8*/	5,24,1,3,34,2,1,119,2,6,26,1,3,26,2,2,
/* out0177_em-eta17-phi8*/	5,24,0,4,24,1,1,112,1,1,119,2,4,26,2,3,
/* out0178_em-eta18-phi8*/	5,23,0,1,24,0,3,112,1,4,15,1,2,26,2,1,
/* out0179_em-eta19-phi8*/	1,24,0,1,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	2,95,1,6,96,0,2,
/* out0185_em-eta5-phi9*/	12,91,1,2,91,2,2,92,0,5,92,1,9,99,0,12,99,1,13,99,2,14,85,1,3,86,0,5,95,0,3,95,1,8,95,2,15,
/* out0186_em-eta6-phi9*/	8,81,1,12,91,2,10,92,0,6,74,0,2,74,1,1,85,1,11,85,2,8,86,0,5,
/* out0187_em-eta7-phi9*/	9,70,1,3,80,2,3,81,0,16,81,1,2,81,2,1,73,1,5,74,0,13,74,2,1,85,2,2,
/* out0188_em-eta8-phi9*/	8,70,0,4,70,1,10,70,2,6,62,0,7,62,1,5,73,1,1,73,2,3,74,2,2,
/* out0189_em-eta9-phi9*/	7,58,1,5,58,2,2,59,0,1,70,0,6,70,2,3,62,0,7,62,2,7,
/* out0190_em-eta10-phi9*/	5,58,0,1,58,1,2,58,2,11,50,0,3,50,1,9,
/* out0191_em-eta11-phi9*/	12,46,1,1,46,2,1,47,0,2,47,1,3,58,0,2,58,2,2,135,1,7,135,2,6,136,0,1,50,0,1,50,1,1,50,2,9,
/* out0192_em-eta12-phi9*/	8,46,2,7,47,0,3,128,1,1,135,0,2,135,2,9,38,1,6,39,0,1,50,2,2,
/* out0193_em-eta13-phi9*/	9,35,1,6,46,2,2,127,1,1,127,2,4,128,0,4,128,1,1,135,0,1,38,1,4,38,2,3,
/* out0194_em-eta14-phi9*/	7,35,0,6,35,1,1,120,1,2,127,2,6,128,0,1,27,0,2,38,2,4,
/* out0195_em-eta15-phi9*/	7,24,1,2,34,2,1,35,0,3,120,0,2,120,1,5,26,1,2,27,0,3,
/* out0196_em-eta16-phi9*/	4,24,1,5,120,0,6,26,1,2,27,0,1,
/* out0197_em-eta17-phi9*/	7,24,0,2,24,1,1,112,1,2,112,2,3,120,0,1,15,1,3,26,2,1,
/* out0198_em-eta18-phi9*/	4,24,0,3,112,1,5,112,2,1,15,1,4,
/* out0199_em-eta19-phi9*/	1,24,0,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	2,96,0,10,96,2,1,
/* out0205_em-eta5-phi10*/	10,92,0,1,92,1,7,92,2,11,93,0,8,93,2,1,86,0,4,86,1,14,87,0,1,96,0,4,96,2,13,
/* out0206_em-eta6-phi10*/	11,81,1,2,81,2,4,82,0,6,82,1,8,92,0,4,92,2,5,74,1,5,75,0,3,86,0,2,86,1,1,86,2,15,
/* out0207_em-eta7-phi10*/	8,71,1,10,81,2,11,82,0,3,63,0,1,74,0,1,74,1,10,74,2,9,75,0,1,
/* out0208_em-eta8-phi10*/	6,59,1,2,70,2,6,71,0,12,62,1,8,63,0,7,74,2,4,
/* out0209_em-eta9-phi10*/	7,59,0,4,59,1,11,70,2,1,51,0,4,62,1,3,62,2,8,63,0,1,
/* out0210_em-eta10-phi10*/	6,47,1,4,58,2,1,59,0,9,50,1,4,51,0,8,62,2,1,
/* out0211_em-eta11-phi10*/	10,47,0,2,47,1,8,47,2,1,136,0,11,136,2,2,39,0,3,39,1,1,50,1,2,50,2,3,51,2,1,
/* out0212_em-eta12-phi10*/	8,35,1,1,47,0,8,47,2,1,128,1,9,135,2,1,136,0,1,136,2,4,39,0,9,
/* out0213_em-eta13-phi10*/	10,35,1,7,35,2,1,128,0,5,128,1,3,128,2,2,27,1,1,38,1,1,38,2,1,39,0,2,39,2,2,
/* out0214_em-eta14-phi10*/	7,35,0,2,35,1,1,35,2,3,120,1,4,128,0,5,27,0,4,27,1,2,
/* out0215_em-eta15-phi10*/	7,24,1,1,35,0,4,35,2,1,120,1,5,120,2,3,27,0,5,27,2,1,
/* out0216_em-eta16-phi10*/	6,24,1,3,24,2,2,120,0,4,120,2,2,27,0,1,27,2,3,
/* out0217_em-eta17-phi10*/	5,24,2,4,112,2,4,120,0,2,15,1,1,15,2,4,
/* out0218_em-eta18-phi10*/	6,24,0,1,24,2,3,112,1,2,112,2,4,15,1,3,15,2,1,
/* out0219_em-eta19-phi10*/	3,24,0,1,24,2,1,112,1,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	3,87,0,1,87,1,3,96,2,1,
/* out0225_em-eta5-phi11*/	8,82,1,1,83,1,4,93,0,8,93,2,15,87,0,14,87,1,9,87,2,9,96,2,1,
/* out0226_em-eta6-phi11*/	11,72,1,1,82,0,3,82,1,7,82,2,14,83,0,4,75,0,9,75,1,12,75,2,2,86,1,1,86,2,1,87,2,3,
/* out0227_em-eta7-phi11*/	10,71,1,6,71,2,6,72,0,4,72,1,3,82,0,4,82,2,2,63,0,1,63,1,7,75,0,3,75,2,10,
/* out0228_em-eta8-phi11*/	8,59,1,1,60,0,1,60,1,4,71,0,4,71,2,10,63,0,6,63,1,5,63,2,7,
/* out0229_em-eta9-phi11*/	6,59,1,2,59,2,11,60,0,3,51,0,1,51,1,9,63,2,5,
/* out0230_em-eta10-phi11*/	9,47,1,1,47,2,1,48,0,1,48,1,4,59,0,2,59,2,5,51,0,3,51,1,3,51,2,7,
/* out0231_em-eta11-phi11*/	7,47,2,8,48,0,3,129,1,2,136,0,3,136,2,7,39,1,7,51,2,4,
/* out0232_em-eta12-phi11*/	11,36,1,4,47,0,1,47,2,5,128,1,2,128,2,3,129,0,3,129,1,2,136,2,3,39,0,1,39,1,4,39,2,4,
/* out0233_em-eta13-phi11*/	7,35,2,3,36,0,4,121,1,1,128,2,9,129,0,1,27,1,1,39,2,6,
/* out0234_em-eta14-phi11*/	8,25,1,1,35,2,6,120,2,1,121,0,2,121,1,3,128,0,1,128,2,2,27,1,6,
/* out0235_em-eta15-phi11*/	7,25,0,1,25,1,3,35,2,2,120,2,5,121,0,2,27,1,2,27,2,3,
/* out0236_em-eta16-phi11*/	5,24,2,2,25,0,3,113,1,2,120,2,4,27,2,4,
/* out0237_em-eta17-phi11*/	7,24,2,3,112,2,1,113,0,2,113,1,2,120,2,1,15,2,4,27,2,1,
/* out0238_em-eta18-phi11*/	6,14,1,2,24,2,1,112,2,3,113,0,2,15,1,1,15,2,3,
/* out0239_em-eta19-phi11*/	3,14,1,3,112,1,1,15,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	1,88,0,7,
/* out0245_em-eta5-phi12*/	9,83,1,12,83,2,8,84,0,3,76,0,5,76,1,7,87,1,4,87,2,4,88,0,8,88,2,8,
/* out0246_em-eta6-phi12*/	12,72,1,7,72,2,3,73,0,1,73,1,1,83,0,12,83,2,6,64,1,2,75,1,4,75,2,1,76,0,11,76,1,1,76,2,7,
/* out0247_em-eta7-phi12*/	8,72,0,10,72,1,5,72,2,9,63,1,1,64,0,14,64,1,4,64,2,1,75,2,3,
/* out0248_em-eta8-phi12*/	10,60,0,1,60,1,12,60,2,5,72,0,2,52,0,4,52,1,3,63,1,3,63,2,4,64,0,2,64,2,3,
/* out0249_em-eta9-phi12*/	6,48,1,3,60,0,11,60,2,2,51,1,2,52,0,11,52,2,1,
/* out0250_em-eta10-phi12*/	9,48,0,2,48,1,9,48,2,3,40,0,4,40,1,1,51,1,2,51,2,4,52,0,1,52,2,1,
/* out0251_em-eta11-phi12*/	7,36,1,2,48,0,9,48,2,1,129,1,8,129,2,1,39,1,1,40,0,9,
/* out0252_em-eta12-phi12*/	10,36,1,9,36,2,1,129,0,6,129,1,4,129,2,3,28,0,1,39,1,3,39,2,2,40,0,1,40,2,1,
/* out0253_em-eta13-phi12*/	6,36,0,7,36,2,1,121,1,6,129,0,5,28,0,6,39,2,2,
/* out0254_em-eta14-phi12*/	7,25,1,4,36,0,3,121,0,3,121,1,5,121,2,1,27,1,2,28,0,4,
/* out0255_em-eta15-phi12*/	6,25,0,1,25,1,5,121,0,7,16,0,1,27,1,2,27,2,2,
/* out0256_em-eta16-phi12*/	4,25,0,5,113,1,6,16,0,3,27,2,2,
/* out0257_em-eta17-phi12*/	6,14,2,2,25,0,2,113,0,3,113,1,3,15,2,1,16,0,3,
/* out0258_em-eta18-phi12*/	4,14,1,3,14,2,1,113,0,4,15,2,3,
/* out0259_em-eta19-phi12*/	3,14,1,3,113,0,1,15,1,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	4,77,0,1,77,1,4,88,0,1,88,2,3,
/* out0265_em-eta5-phi13*/	11,73,1,3,73,2,1,74,0,1,83,2,1,84,0,13,84,2,14,76,1,7,77,0,15,77,1,3,77,2,4,88,2,5,
/* out0266_em-eta6-phi13*/	9,73,0,10,73,1,12,73,2,6,83,2,1,64,1,2,65,0,12,65,1,2,76,1,1,76,2,9,
/* out0267_em-eta7-phi13*/	8,61,1,15,61,2,1,72,2,4,73,0,5,53,0,3,64,1,8,64,2,8,65,0,3,
/* out0268_em-eta8-phi13*/	6,49,1,2,60,2,5,61,0,13,52,1,9,53,0,5,64,2,4,
/* out0269_em-eta9-phi13*/	5,49,0,4,49,1,9,60,2,4,52,1,4,52,2,11,
/* out0270_em-eta10-phi13*/	6,37,1,1,48,2,8,49,0,4,40,1,10,41,0,1,52,2,2,
/* out0271_em-eta11-phi13*/	10,36,1,1,37,0,2,37,1,5,48,0,1,48,2,4,129,2,3,130,0,9,40,0,2,40,1,2,40,2,6,
/* out0272_em-eta12-phi13*/	7,36,2,7,37,0,2,122,1,3,129,2,8,130,0,1,28,1,5,40,2,4,
/* out0273_em-eta13-phi13*/	12,26,1,1,36,0,1,36,2,7,121,1,1,121,2,2,122,0,3,122,1,2,129,0,1,129,2,1,28,0,3,28,1,4,28,2,1,
/* out0274_em-eta14-phi13*/	7,25,1,2,25,2,2,26,0,1,36,0,1,121,2,9,28,0,2,28,2,4,
/* out0275_em-eta15-phi13*/	8,25,1,1,25,2,5,114,1,1,121,0,2,121,2,3,16,0,1,16,1,3,28,2,1,
/* out0276_em-eta16-phi13*/	6,25,0,2,25,2,3,113,1,3,113,2,4,16,0,3,16,1,1,
/* out0277_em-eta17-phi13*/	4,14,2,3,25,0,2,113,2,5,16,0,3,
/* out0278_em-eta18-phi13*/	5,14,2,4,113,0,3,113,2,1,16,0,2,16,2,1,
/* out0279_em-eta19-phi13*/	2,14,1,2,113,0,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	4,77,1,4,78,0,12,78,1,6,78,2,7,
/* out0285_em-eta5-phi14*/	12,74,0,15,74,1,10,74,2,7,84,2,2,65,1,1,66,0,10,66,1,2,77,1,5,77,2,12,78,0,2,78,1,7,78,2,5,
/* out0286_em-eta6-phi14*/	8,62,1,12,73,2,9,74,2,8,54,0,1,65,0,1,65,1,13,65,2,9,66,0,3,
/* out0287_em-eta7-phi14*/	9,50,1,1,61,1,1,61,2,10,62,0,10,62,1,1,53,0,1,53,1,12,54,0,2,65,2,7,
/* out0288_em-eta8-phi14*/	9,49,1,2,49,2,1,50,0,3,50,1,5,61,0,3,61,2,5,53,0,7,53,1,1,53,2,10,
/* out0289_em-eta9-phi14*/	7,49,0,2,49,1,3,49,2,11,41,0,7,41,1,7,52,2,1,53,2,1,
/* out0290_em-eta10-phi14*/	7,37,1,5,37,2,1,49,0,6,49,2,2,40,1,2,41,0,8,41,2,3,
/* out0291_em-eta11-phi14*/	9,37,0,3,37,1,5,37,2,3,130,0,6,130,2,12,29,0,4,29,1,1,40,1,1,40,2,4,
/* out0292_em-eta12-phi14*/	8,26,1,2,37,0,7,122,1,9,122,2,2,130,2,2,28,1,3,29,0,5,40,2,1,
/* out0293_em-eta13-phi14*/	6,26,1,8,122,0,8,122,1,2,122,2,2,28,1,4,28,2,3,
/* out0294_em-eta14-phi14*/	6,26,0,6,26,1,1,114,1,5,121,2,1,122,0,3,28,2,6,
/* out0295_em-eta15-phi14*/	7,15,1,1,25,2,3,26,0,1,114,0,2,114,1,6,16,1,4,28,2,1,
/* out0296_em-eta16-phi14*/	6,15,1,2,25,2,2,113,2,1,114,0,5,16,1,4,16,2,1,
/* out0297_em-eta17-phi14*/	7,14,2,1,15,0,2,15,1,1,25,2,1,107,1,1,113,2,3,16,2,3,
/* out0298_em-eta18-phi14*/	4,14,2,4,107,1,2,113,2,2,16,2,3,
/* out0299_em-eta19-phi14*/	2,14,1,2,107,1,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	3,67,1,9,78,0,2,78,2,2,
/* out0305_em-eta5-phi15*/	11,63,1,13,74,1,5,55,0,1,66,0,2,66,1,14,66,2,9,67,0,16,67,1,1,67,2,1,78,1,3,78,2,2,
/* out0306_em-eta6-phi15*/	12,51,1,2,62,1,3,62,2,11,63,0,10,63,1,2,74,1,1,74,2,1,54,0,4,54,1,13,55,0,1,66,0,1,66,2,7,
/* out0307_em-eta7-phi15*/	10,50,1,5,50,2,3,51,0,2,51,1,3,62,0,6,62,2,5,42,1,2,53,1,3,54,0,9,54,2,8,
/* out0308_em-eta8-phi15*/	6,50,0,8,50,1,5,50,2,7,42,0,10,42,1,2,53,2,5,
/* out0309_em-eta9-phi15*/	6,38,1,10,49,2,2,50,0,5,41,1,9,41,2,3,42,0,3,
/* out0310_em-eta10-phi15*/	6,37,2,2,38,0,8,38,1,4,29,1,2,30,0,1,41,2,10,
/* out0311_em-eta11-phi15*/	9,27,1,2,37,2,8,38,0,1,123,0,16,123,1,4,123,2,2,130,2,2,29,0,2,29,1,9,
/* out0312_em-eta12-phi15*/	11,26,1,2,26,2,2,27,0,1,27,1,2,37,0,2,37,2,2,115,1,1,122,2,6,123,2,8,29,0,4,29,2,5,
/* out0313_em-eta13-phi15*/	9,26,1,2,26,2,5,115,1,3,122,0,1,122,2,6,17,0,2,17,1,3,29,0,1,29,2,2,
/* out0314_em-eta14-phi15*/	7,26,0,5,26,2,2,114,1,3,114,2,4,115,0,1,122,0,1,17,0,6,
/* out0315_em-eta15-phi15*/	7,15,1,4,26,0,2,114,0,2,114,1,1,114,2,5,16,1,1,17,0,4,
/* out0316_em-eta16-phi15*/	4,15,1,5,114,0,6,16,1,3,16,2,2,
/* out0317_em-eta17-phi15*/	4,15,0,3,107,1,1,107,2,4,16,2,4,
/* out0318_em-eta18-phi15*/	4,14,2,1,15,0,3,107,1,4,16,2,2,
/* out0319_em-eta19-phi15*/	2,14,1,1,107,1,2,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	3,56,1,2,67,1,6,67,2,2,
/* out0325_em-eta5-phi16*/	12,52,1,4,63,1,1,63,2,12,64,0,15,64,1,14,64,2,12,55,0,5,55,1,14,55,2,2,56,0,5,56,1,4,67,2,13,
/* out0326_em-eta6-phi16*/	12,51,1,7,51,2,5,52,0,3,52,1,4,63,0,6,63,2,4,43,0,1,43,1,4,54,1,3,54,2,2,55,0,9,55,2,8,
/* out0327_em-eta7-phi16*/	7,39,1,1,51,0,13,51,1,4,51,2,6,42,1,4,43,0,11,54,2,6,
/* out0328_em-eta8-phi16*/	6,39,0,2,39,1,12,50,2,6,42,0,2,42,1,8,42,2,9,
/* out0329_em-eta9-phi16*/	7,38,1,2,38,2,10,39,0,5,30,0,2,30,1,7,42,0,1,42,2,6,
/* out0330_em-eta10-phi16*/	6,27,1,1,38,0,7,38,2,6,30,0,11,30,1,1,30,2,1,
/* out0331_em-eta11-phi16*/	8,27,1,10,27,2,1,123,1,10,18,0,1,29,1,4,29,2,3,30,0,2,30,2,1,
/* out0332_em-eta12-phi16*/	8,27,0,8,27,1,1,115,1,5,115,2,1,123,1,2,123,2,6,18,0,2,29,2,6,
/* out0333_em-eta13-phi16*/	7,16,1,2,26,2,4,27,0,2,115,0,2,115,1,7,115,2,1,17,1,7,
/* out0334_em-eta14-phi16*/	8,16,1,3,26,0,1,26,2,3,114,2,1,115,0,7,17,0,2,17,1,2,17,2,2,
/* out0335_em-eta15-phi16*/	7,15,1,2,15,2,3,16,0,1,108,1,3,114,2,5,17,0,2,17,2,3,
/* out0336_em-eta16-phi16*/	10,15,1,1,15,2,3,107,2,2,108,0,1,108,1,2,114,0,1,114,2,1,7,1,1,7,2,1,17,2,1,
/* out0337_em-eta17-phi16*/	3,15,0,3,107,2,6,7,1,3,
/* out0338_em-eta18-phi16*/	5,15,0,3,107,0,2,107,1,2,107,2,1,7,1,2,
/* out0339_em-eta19-phi16*/	1,107,1,2,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	1,56,1,4,
/* out0345_em-eta5-phi17*/	15,52,1,6,52,2,9,53,0,12,53,1,8,53,2,4,64,0,1,64,1,2,64,2,4,44,0,4,44,1,8,55,1,2,55,2,3,56,0,11,56,1,6,56,2,16,
/* out0346_em-eta6-phi17*/	9,40,1,6,51,2,1,52,0,13,52,1,2,52,2,7,43,1,10,43,2,1,44,0,12,55,2,3,
/* out0347_em-eta7-phi17*/	10,39,1,1,39,2,1,40,0,7,40,1,10,51,0,1,51,2,4,31,1,1,43,0,3,43,1,2,43,2,15,
/* out0348_em-eta8-phi17*/	8,39,0,2,39,1,2,39,2,14,40,0,1,31,0,9,31,1,7,42,2,1,43,0,1,
/* out0349_em-eta9-phi17*/	6,28,1,9,39,0,7,39,2,1,30,1,7,30,2,1,31,0,7,
/* out0350_em-eta10-phi17*/	4,28,0,6,28,1,7,30,1,1,30,2,11,
/* out0351_em-eta11-phi17*/	7,27,2,10,28,0,2,116,0,12,116,1,5,18,0,1,18,1,7,30,2,2,
/* out0352_em-eta12-phi17*/	7,27,0,4,27,2,5,115,2,3,116,0,4,116,2,8,18,0,8,18,1,1,
/* out0353_em-eta13-phi17*/	6,16,1,7,27,0,1,115,0,1,115,2,10,17,1,4,18,0,4,
/* out0354_em-eta14-phi17*/	6,16,0,3,16,1,4,108,1,3,115,0,5,115,2,1,17,2,6,
/* out0355_em-eta15-phi17*/	5,15,2,2,16,0,4,108,1,7,7,2,1,17,2,4,
/* out0356_em-eta16-phi17*/	4,15,2,5,108,0,5,108,1,1,7,2,5,
/* out0357_em-eta17-phi17*/	6,15,0,1,15,2,3,107,0,1,107,2,3,108,0,2,7,1,3,
/* out0358_em-eta18-phi17*/	3,15,0,1,107,0,10,7,1,2,
/* out0359_em-eta19-phi17*/	2,107,0,3,107,1,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	1,45,1,5,
/* out0365_em-eta5-phi18*/	15,41,1,9,41,2,6,42,0,4,42,1,2,42,2,1,53,0,4,53,1,8,53,2,12,33,0,3,33,1,2,44,1,8,44,2,4,45,0,16,45,1,10,45,2,9,
/* out0366_em-eta6-phi18*/	9,30,1,1,40,2,6,41,0,13,41,1,7,41,2,2,32,0,1,32,1,10,33,0,3,44,2,12,
/* out0367_em-eta7-phi18*/	10,29,1,1,29,2,1,30,0,1,30,1,4,40,0,7,40,2,10,31,1,1,32,0,15,32,1,2,32,2,3,
/* out0368_em-eta8-phi18*/	8,29,0,2,29,1,14,29,2,2,40,0,1,20,0,1,31,1,7,31,2,9,32,2,1,
/* out0369_em-eta9-phi18*/	6,28,2,9,29,0,7,29,1,1,19,0,1,19,1,7,31,2,7,
/* out0370_em-eta10-phi18*/	4,28,0,6,28,2,7,19,0,11,19,1,1,
/* out0371_em-eta11-phi18*/	7,17,1,10,28,0,2,110,0,1,116,1,9,18,1,7,18,2,1,19,0,2,
/* out0372_em-eta12-phi18*/	7,17,0,4,17,1,5,109,1,3,116,1,2,116,2,8,18,1,1,18,2,8,
/* out0373_em-eta13-phi18*/	6,16,2,7,17,0,1,109,0,1,109,1,10,8,1,4,18,2,4,
/* out0374_em-eta14-phi18*/	6,16,0,3,16,2,4,108,2,3,109,0,5,109,1,1,8,0,6,
/* out0375_em-eta15-phi18*/	5,7,1,2,16,0,4,108,2,7,7,2,1,8,0,4,
/* out0376_em-eta16-phi18*/	4,7,1,5,108,0,5,108,2,1,7,2,5,
/* out0377_em-eta17-phi18*/	8,7,0,1,7,1,3,103,1,1,103,2,3,108,0,2,7,0,3,7,1,2,7,2,1,
/* out0378_em-eta18-phi18*/	3,7,0,1,103,1,4,7,1,2,
/* out0379_em-eta19-phi18*/	1,103,1,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	3,34,1,8,45,1,1,45,2,1,
/* out0385_em-eta5-phi19*/	13,31,1,12,31,2,1,41,2,4,42,0,12,42,1,14,42,2,15,33,0,2,33,1,14,33,2,5,34,0,16,34,1,5,34,2,2,45,2,6,
/* out0386_em-eta6-phi19*/	12,30,1,5,30,2,7,31,0,6,31,1,4,41,0,3,41,2,4,21,0,2,21,1,3,32,1,4,32,2,1,33,0,8,33,2,9,
/* out0387_em-eta7-phi19*/	7,29,2,1,30,0,13,30,1,6,30,2,4,20,1,4,21,0,6,32,2,11,
/* out0388_em-eta8-phi19*/	6,19,1,6,29,0,2,29,2,12,20,0,9,20,1,8,20,2,2,
/* out0389_em-eta9-phi19*/	7,18,1,10,18,2,2,29,0,5,19,1,7,19,2,2,20,0,6,20,2,1,
/* out0390_em-eta10-phi19*/	6,17,2,1,18,0,7,18,1,6,19,0,1,19,1,1,19,2,11,
/* out0391_em-eta11-phi19*/	10,17,1,1,17,2,10,110,0,12,110,1,5,110,2,1,9,0,3,9,1,4,18,2,1,19,0,1,19,2,2,
/* out0392_em-eta12-phi19*/	8,17,0,8,17,2,1,109,1,1,109,2,5,110,0,3,110,2,7,9,0,6,18,2,2,
/* out0393_em-eta13-phi19*/	7,8,1,4,16,2,2,17,0,2,109,0,2,109,1,1,109,2,7,8,1,7,
/* out0394_em-eta14-phi19*/	8,8,0,1,8,1,3,16,2,3,104,1,1,109,0,7,8,0,2,8,1,2,8,2,2,
/* out0395_em-eta15-phi19*/	7,7,1,3,7,2,2,16,0,1,104,1,5,108,2,3,8,0,3,8,2,2,
/* out0396_em-eta16-phi19*/	10,7,1,3,7,2,1,103,2,2,104,0,1,104,1,1,108,0,1,108,2,2,7,0,3,7,2,2,8,0,1,
/* out0397_em-eta17-phi19*/	3,7,0,3,103,2,6,7,0,8,
/* out0398_em-eta18-phi19*/	5,7,0,3,103,1,3,103,2,1,7,0,1,7,1,1,
/* out0399_em-eta19-phi19*/	1,103,1,2,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	4,23,0,2,23,2,2,34,1,3,34,2,6,
/* out0405_em-eta5-phi20*/	10,21,0,11,21,1,2,31,2,13,22,0,9,22,1,14,22,2,2,23,0,2,23,1,3,33,2,1,34,2,8,
/* out0406_em-eta6-phi20*/	12,20,1,11,20,2,3,21,0,2,21,2,1,30,2,2,31,0,10,31,2,2,21,1,13,21,2,4,22,0,7,22,2,1,33,2,1,
/* out0407_em-eta7-phi20*/	10,19,1,3,19,2,5,20,0,6,20,1,5,30,0,2,30,2,3,11,1,3,20,1,2,21,0,8,21,2,9,
/* out0408_em-eta8-phi20*/	6,19,0,8,19,1,7,19,2,5,11,0,5,20,1,2,20,2,10,
/* out0409_em-eta9-phi20*/	6,10,1,2,18,2,10,19,0,5,10,0,3,10,1,9,20,2,3,
/* out0410_em-eta10-phi20*/	6,9,1,2,18,0,8,18,2,4,9,1,2,10,0,10,19,2,1,
/* out0411_em-eta11-phi20*/	8,9,1,8,17,2,2,18,0,1,106,0,2,110,1,11,110,2,1,9,1,9,9,2,2,
/* out0412_em-eta12-phi20*/	11,8,1,2,8,2,2,9,0,2,9,1,2,17,0,1,17,2,2,105,1,6,109,2,1,110,2,7,9,0,5,9,2,4,
/* out0413_em-eta13-phi20*/	9,8,1,5,8,2,2,105,0,1,105,1,6,109,2,3,8,1,3,8,2,2,9,0,2,9,2,1,
/* out0414_em-eta14-phi20*/	7,8,0,5,8,1,2,104,1,4,104,2,3,105,0,1,109,0,1,8,2,6,
/* out0415_em-eta15-phi20*/	7,7,2,4,8,0,2,104,0,2,104,1,5,104,2,1,0,1,1,8,2,4,
/* out0416_em-eta16-phi20*/	4,7,2,5,104,0,6,0,0,2,0,1,3,
/* out0417_em-eta17-phi20*/	4,7,0,3,103,0,2,103,2,4,0,0,4,
/* out0418_em-eta18-phi20*/	6,0,1,1,7,0,3,103,0,5,103,1,2,0,0,2,7,0,1,
/* out0419_em-eta19-phi20*/	2,0,1,1,103,1,1,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	4,13,1,4,23,0,7,23,1,6,23,2,12,
/* out0425_em-eta5-phi21*/	12,13,0,2,21,0,3,21,1,14,21,2,7,12,1,1,13,0,12,13,1,5,22,1,2,22,2,10,23,0,5,23,1,7,23,2,2,
/* out0426_em-eta6-phi21*/	8,12,1,9,20,2,12,21,2,8,12,0,9,12,1,13,12,2,1,21,2,1,22,2,3,
/* out0427_em-eta7-phi21*/	9,11,1,10,11,2,1,19,2,1,20,0,10,20,2,1,11,1,12,11,2,1,12,0,7,21,2,2,
/* out0428_em-eta8-phi21*/	9,10,1,1,10,2,2,11,0,3,11,1,5,19,0,3,19,2,5,11,0,10,11,1,1,11,2,7,
/* out0429_em-eta9-phi21*/	7,10,0,2,10,1,11,10,2,3,3,0,1,10,1,7,10,2,7,11,0,1,
/* out0430_em-eta10-phi21*/	7,9,1,1,9,2,5,10,0,6,10,1,2,2,1,2,10,0,3,10,2,8,
/* out0431_em-eta11-phi21*/	9,9,0,3,9,1,3,9,2,5,106,0,12,106,2,6,2,0,4,2,1,1,9,1,1,9,2,4,
/* out0432_em-eta12-phi21*/	8,8,2,2,9,0,7,105,1,2,105,2,9,106,2,2,1,1,3,2,0,1,9,2,5,
/* out0433_em-eta13-phi21*/	6,8,2,8,105,0,8,105,1,2,105,2,2,1,0,3,1,1,4,
/* out0434_em-eta14-phi21*/	6,8,0,6,8,2,1,101,1,1,104,2,5,105,0,3,1,0,6,
/* out0435_em-eta15-phi21*/	7,1,1,3,7,2,1,8,0,1,104,0,2,104,2,6,0,1,4,1,0,1,
/* out0436_em-eta16-phi21*/	6,1,1,2,7,2,2,100,1,1,104,0,5,0,0,1,0,1,4,
/* out0437_em-eta17-phi21*/	9,0,1,1,0,2,1,1,0,1,1,1,1,7,0,2,7,2,1,100,1,3,103,0,3,0,0,3,
/* out0438_em-eta18-phi21*/	4,0,1,4,100,1,2,103,0,6,0,0,3,
/* out0439_em-eta19-phi21*/	3,0,1,2,100,0,1,103,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	3,6,0,4,13,1,4,13,2,1,
/* out0445_em-eta5-phi22*/	11,6,1,1,12,1,1,12,2,3,13,0,14,13,2,14,5,1,7,6,0,5,6,2,1,13,0,4,13,1,3,13,2,15,
/* out0446_em-eta6-phi22*/	9,6,1,1,12,0,10,12,1,6,12,2,12,4,1,2,5,0,9,5,1,1,12,1,2,12,2,12,
/* out0447_em-eta7-phi22*/	8,5,1,4,11,1,1,11,2,15,12,0,5,4,0,8,4,1,8,11,2,3,12,2,3,
/* out0448_em-eta8-phi22*/	6,4,1,5,10,2,2,11,0,13,3,1,9,4,0,4,11,2,5,
/* out0449_em-eta9-phi22*/	7,3,2,1,4,0,1,4,1,4,10,0,4,10,2,9,3,0,11,3,1,4,
/* out0450_em-eta10-phi22*/	6,3,1,8,9,2,1,10,0,4,2,1,10,3,0,2,10,2,1,
/* out0451_em-eta11-phi22*/	12,2,2,1,3,0,1,3,1,4,9,0,2,9,2,5,102,1,3,102,2,3,106,0,2,106,2,7,2,0,6,2,1,2,2,2,2,
/* out0452_em-eta12-phi22*/	9,2,1,7,2,2,1,9,0,2,102,0,3,102,1,8,105,2,3,106,2,1,1,1,5,2,0,4,
/* out0453_em-eta13-phi22*/	12,2,0,1,2,1,7,8,2,1,101,1,2,101,2,2,102,0,1,102,1,1,105,0,3,105,2,2,1,0,1,1,1,4,1,2,3,
/* out0454_em-eta14-phi22*/	8,1,1,2,1,2,3,2,0,4,8,0,1,101,1,9,101,2,2,1,0,4,1,2,2,
/* out0455_em-eta15-phi22*/	10,1,0,1,1,1,5,1,2,1,100,2,1,101,0,5,101,1,3,104,2,1,0,1,3,0,2,1,1,0,1,
/* out0456_em-eta16-phi22*/	6,1,0,2,1,1,3,100,1,4,100,2,3,0,1,1,0,2,3,
/* out0457_em-eta17-phi22*/	6,0,2,3,1,0,3,100,0,1,100,1,5,100,2,1,0,2,3,
/* out0458_em-eta18-phi22*/	6,0,1,2,0,2,3,100,0,4,100,1,1,0,0,1,0,2,2,
/* out0459_em-eta19-phi22*/	3,0,1,3,0,2,1,100,0,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	2,6,0,5,6,2,1,
/* out0465_em-eta5-phi23*/	8,6,0,4,6,1,8,6,2,16,13,2,2,5,1,7,5,2,5,6,0,2,6,2,14,
/* out0466_em-eta6-phi23*/	10,5,1,3,5,2,11,6,0,12,6,1,6,12,0,1,12,2,1,4,1,2,5,0,7,5,1,1,5,2,11,
/* out0467_em-eta7-phi23*/	6,5,0,14,5,1,9,5,2,5,4,0,1,4,1,4,4,2,14,
/* out0468_em-eta8-phi23*/	8,4,0,1,4,1,5,4,2,16,5,0,2,3,1,3,3,2,4,4,0,3,4,2,2,
/* out0469_em-eta9-phi23*/	5,3,2,6,4,0,14,4,1,2,3,0,1,3,2,11,
/* out0470_em-eta10-phi23*/	7,3,0,2,3,1,3,3,2,9,2,1,1,2,2,4,3,0,1,3,2,1,
/* out0471_em-eta11-phi23*/	6,2,2,2,3,0,13,3,1,1,102,1,1,102,2,9,2,2,9,
/* out0472_em-eta12-phi23*/	8,2,1,1,2,2,9,102,0,7,102,1,3,102,2,4,1,2,1,2,0,1,2,2,1,
/* out0473_em-eta13-phi23*/	6,2,0,8,2,1,1,2,2,3,101,2,6,102,0,5,1,2,6,
/* out0474_em-eta14-phi23*/	6,1,2,7,2,0,3,101,0,3,101,1,1,101,2,6,1,2,4,
/* out0475_em-eta15-phi23*/	5,1,0,1,1,2,5,100,2,1,101,0,8,0,2,1,
/* out0476_em-eta16-phi23*/	3,1,0,5,100,2,7,0,2,3,
/* out0477_em-eta17-phi23*/	5,0,2,2,1,0,3,100,0,3,100,2,3,0,2,3,
/* out0478_em-eta18-phi23*/	2,0,2,5,100,0,5,
/* out0479_em-eta19-phi23*/	3,0,1,2,0,2,1,100,0,1
};