parameter integer matrixH [0:4212] = {
/* num inputs = 133(in0-in132) */
/* num outputs = 560(out0-out559) */
//* max inputs per outputs = 11 */
//* total number of input in adders 1244 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	0, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	0, 
/* out0033_had-eta13-phi1*/	0, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	0, 
/* out0036_had-eta16-phi1*/	0, 
/* out0037_had-eta17-phi1*/	0, 
/* out0038_had-eta18-phi1*/	0, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	0, 
/* out0045_had-eta5-phi2*/	0, 
/* out0046_had-eta6-phi2*/	0, 
/* out0047_had-eta7-phi2*/	0, 
/* out0048_had-eta8-phi2*/	0, 
/* out0049_had-eta9-phi2*/	0, 
/* out0050_had-eta10-phi2*/	0, 
/* out0051_had-eta11-phi2*/	1, 104, 2, 3, 
/* out0052_had-eta12-phi2*/	2, 104, 1, 4, 104, 2, 1, 
/* out0053_had-eta13-phi2*/	1, 103, 2, 2, 
/* out0054_had-eta14-phi2*/	2, 103, 1, 3, 103, 2, 2, 
/* out0055_had-eta15-phi2*/	1, 103, 1, 1, 
/* out0056_had-eta16-phi2*/	1, 102, 2, 3, 
/* out0057_had-eta17-phi2*/	2, 102, 1, 3, 102, 2, 1, 
/* out0058_had-eta18-phi2*/	1, 102, 1, 1, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 110, 0, 10, 
/* out0062_had-eta2-phi3*/	2, 110, 0, 6, 110, 1, 11, 
/* out0063_had-eta3-phi3*/	2, 109, 0, 13, 110, 1, 5, 
/* out0064_had-eta4-phi3*/	2, 109, 0, 3, 109, 1, 14, 
/* out0065_had-eta5-phi3*/	1, 109, 1, 2, 
/* out0066_had-eta6-phi3*/	2, 63, 0, 1, 63, 1, 1, 
/* out0067_had-eta7-phi3*/	3, 62, 2, 5, 63, 0, 1, 63, 1, 13, 
/* out0068_had-eta8-phi3*/	2, 62, 1, 10, 62, 2, 8, 
/* out0069_had-eta9-phi3*/	2, 61, 2, 9, 62, 1, 2, 
/* out0070_had-eta10-phi3*/	2, 61, 1, 9, 61, 2, 2, 
/* out0071_had-eta11-phi3*/	4, 60, 2, 7, 61, 1, 1, 104, 0, 1, 104, 2, 11, 
/* out0072_had-eta12-phi3*/	5, 60, 1, 6, 60, 2, 2, 104, 0, 2, 104, 1, 10, 104, 2, 1, 
/* out0073_had-eta13-phi3*/	4, 59, 2, 2, 60, 1, 1, 103, 2, 8, 104, 1, 2, 
/* out0074_had-eta14-phi3*/	5, 59, 1, 2, 59, 2, 4, 103, 0, 1, 103, 1, 5, 103, 2, 3, 
/* out0075_had-eta15-phi3*/	3, 59, 1, 3, 102, 2, 2, 103, 1, 5, 
/* out0076_had-eta16-phi3*/	2, 58, 1, 1, 102, 2, 6, 
/* out0077_had-eta17-phi3*/	3, 58, 1, 3, 102, 1, 4, 102, 2, 1, 
/* out0078_had-eta18-phi3*/	1, 102, 1, 4, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 110, 3, 10, 
/* out0082_had-eta2-phi4*/	2, 110, 2, 11, 110, 3, 6, 
/* out0083_had-eta3-phi4*/	2, 109, 3, 13, 110, 2, 5, 
/* out0084_had-eta4-phi4*/	2, 109, 2, 14, 109, 3, 3, 
/* out0085_had-eta5-phi4*/	1, 109, 2, 2, 
/* out0086_had-eta6-phi4*/	2, 57, 2, 2, 63, 0, 3, 
/* out0087_had-eta7-phi4*/	6, 57, 1, 6, 57, 2, 8, 62, 0, 3, 62, 2, 2, 63, 0, 11, 63, 1, 2, 
/* out0088_had-eta8-phi4*/	5, 56, 2, 4, 57, 1, 2, 62, 0, 13, 62, 1, 2, 62, 2, 1, 
/* out0089_had-eta9-phi4*/	5, 56, 1, 3, 56, 2, 1, 61, 0, 7, 61, 2, 5, 62, 1, 2, 
/* out0090_had-eta10-phi4*/	3, 55, 2, 1, 61, 0, 8, 61, 1, 6, 
/* out0091_had-eta11-phi4*/	4, 60, 0, 5, 60, 2, 7, 100, 1, 8, 104, 0, 6, 
/* out0092_had-eta12-phi4*/	4, 60, 0, 4, 60, 1, 6, 98, 2, 5, 104, 0, 7, 
/* out0093_had-eta13-phi4*/	5, 59, 2, 6, 60, 1, 3, 98, 1, 3, 103, 0, 5, 103, 2, 1, 
/* out0094_had-eta14-phi4*/	4, 59, 0, 1, 59, 1, 2, 59, 2, 3, 103, 0, 8, 
/* out0095_had-eta15-phi4*/	7, 59, 1, 6, 97, 1, 1, 97, 2, 1, 102, 0, 1, 102, 2, 1, 103, 0, 1, 103, 1, 2, 
/* out0096_had-eta16-phi4*/	4, 58, 1, 5, 59, 1, 1, 102, 0, 4, 102, 2, 2, 
/* out0097_had-eta17-phi4*/	3, 58, 1, 3, 102, 0, 4, 102, 1, 1, 
/* out0098_had-eta18-phi4*/	1, 102, 1, 3, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 112, 0, 10, 
/* out0102_had-eta2-phi5*/	2, 112, 0, 6, 112, 1, 11, 
/* out0103_had-eta3-phi5*/	2, 111, 0, 13, 112, 1, 5, 
/* out0104_had-eta4-phi5*/	2, 111, 0, 3, 111, 1, 14, 
/* out0105_had-eta5-phi5*/	1, 111, 1, 2, 
/* out0106_had-eta6-phi5*/	2, 57, 0, 2, 57, 2, 3, 
/* out0107_had-eta7-phi5*/	4, 50, 2, 2, 57, 0, 14, 57, 1, 5, 57, 2, 3, 
/* out0108_had-eta8-phi5*/	4, 50, 1, 1, 56, 0, 6, 56, 2, 11, 57, 1, 3, 
/* out0109_had-eta9-phi5*/	3, 55, 2, 2, 56, 0, 2, 56, 1, 13, 
/* out0110_had-eta10-phi5*/	4, 55, 1, 2, 55, 2, 12, 61, 0, 1, 100, 0, 4, 
/* out0111_had-eta11-phi5*/	6, 54, 2, 1, 55, 1, 9, 60, 0, 3, 98, 2, 2, 100, 0, 9, 100, 1, 8, 
/* out0112_had-eta12-phi5*/	4, 54, 2, 6, 60, 0, 4, 98, 0, 3, 98, 2, 9, 
/* out0113_had-eta13-phi5*/	5, 54, 1, 4, 59, 0, 4, 59, 2, 1, 98, 0, 1, 98, 1, 10, 
/* out0114_had-eta14-phi5*/	4, 59, 0, 7, 97, 2, 8, 98, 1, 1, 103, 0, 1, 
/* out0115_had-eta15-phi5*/	4, 59, 0, 3, 59, 1, 2, 97, 1, 4, 97, 2, 3, 
/* out0116_had-eta16-phi5*/	4, 58, 0, 4, 58, 1, 3, 97, 1, 3, 102, 0, 3, 
/* out0117_had-eta17-phi5*/	4, 58, 0, 4, 58, 1, 1, 96, 2, 2, 102, 0, 3, 
/* out0118_had-eta18-phi5*/	3, 96, 1, 1, 96, 2, 2, 102, 0, 1, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 112, 3, 10, 
/* out0122_had-eta2-phi6*/	2, 112, 2, 11, 112, 3, 6, 
/* out0123_had-eta3-phi6*/	2, 111, 3, 13, 112, 2, 5, 
/* out0124_had-eta4-phi6*/	2, 111, 2, 14, 111, 3, 3, 
/* out0125_had-eta5-phi6*/	1, 111, 2, 2, 
/* out0126_had-eta6-phi6*/	1, 52, 2, 5, 
/* out0127_had-eta7-phi6*/	4, 50, 0, 6, 50, 1, 1, 50, 2, 14, 52, 2, 1, 
/* out0128_had-eta8-phi6*/	3, 49, 2, 4, 50, 1, 13, 56, 0, 4, 
/* out0129_had-eta9-phi6*/	5, 49, 1, 5, 49, 2, 7, 55, 0, 1, 55, 2, 1, 56, 0, 4, 
/* out0130_had-eta10-phi6*/	4, 49, 1, 1, 55, 0, 12, 100, 0, 2, 101, 2, 4, 
/* out0131_had-eta11-phi6*/	8, 48, 2, 1, 54, 0, 1, 54, 2, 3, 55, 0, 3, 55, 1, 5, 100, 0, 1, 101, 1, 6, 101, 2, 11, 
/* out0132_had-eta12-phi6*/	6, 54, 0, 4, 54, 1, 1, 54, 2, 6, 98, 0, 8, 99, 2, 1, 101, 1, 3, 
/* out0133_had-eta13-phi6*/	6, 54, 1, 8, 97, 2, 1, 98, 0, 4, 98, 1, 2, 99, 1, 1, 99, 2, 3, 
/* out0134_had-eta14-phi6*/	5, 53, 2, 6, 54, 1, 1, 59, 0, 1, 97, 0, 5, 97, 2, 3, 
/* out0135_had-eta15-phi6*/	4, 53, 1, 2, 53, 2, 4, 97, 0, 3, 97, 1, 3, 
/* out0136_had-eta16-phi6*/	4, 53, 1, 3, 58, 0, 5, 96, 2, 2, 97, 1, 4, 
/* out0137_had-eta17-phi6*/	2, 58, 0, 3, 96, 2, 5, 
/* out0138_had-eta18-phi6*/	2, 96, 1, 5, 96, 2, 2, 
/* out0139_had-eta19-phi6*/	1, 96, 1, 1, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 114, 0, 10, 
/* out0142_had-eta2-phi7*/	2, 114, 0, 6, 114, 1, 11, 
/* out0143_had-eta3-phi7*/	2, 113, 0, 13, 114, 1, 5, 
/* out0144_had-eta4-phi7*/	2, 113, 0, 3, 113, 1, 14, 
/* out0145_had-eta5-phi7*/	1, 113, 1, 2, 
/* out0146_had-eta6-phi7*/	3, 52, 0, 6, 52, 1, 3, 52, 2, 10, 
/* out0147_had-eta7-phi7*/	3, 50, 0, 7, 51, 2, 7, 52, 1, 12, 
/* out0148_had-eta8-phi7*/	6, 49, 0, 5, 49, 2, 3, 50, 0, 3, 50, 1, 1, 51, 1, 5, 51, 2, 4, 
/* out0149_had-eta9-phi7*/	3, 49, 0, 10, 49, 1, 6, 49, 2, 2, 
/* out0150_had-eta10-phi7*/	3, 48, 2, 11, 49, 1, 4, 101, 0, 2, 
/* out0151_had-eta11-phi7*/	6, 48, 1, 8, 48, 2, 4, 54, 0, 1, 101, 0, 14, 101, 1, 4, 101, 2, 1, 
/* out0152_had-eta12-phi7*/	6, 44, 2, 1, 48, 1, 1, 54, 0, 7, 99, 0, 1, 99, 2, 8, 101, 1, 3, 
/* out0153_had-eta13-phi7*/	8, 44, 2, 1, 53, 0, 1, 53, 2, 1, 54, 0, 3, 54, 1, 2, 99, 0, 1, 99, 1, 5, 99, 2, 4, 
/* out0154_had-eta14-phi7*/	5, 53, 0, 3, 53, 2, 4, 92, 2, 1, 97, 0, 3, 99, 1, 5, 
/* out0155_had-eta15-phi7*/	5, 53, 0, 2, 53, 1, 3, 53, 2, 1, 92, 2, 3, 97, 0, 4, 
/* out0156_had-eta16-phi7*/	7, 53, 1, 5, 92, 1, 1, 92, 2, 1, 96, 0, 2, 96, 2, 2, 97, 0, 1, 97, 1, 1, 
/* out0157_had-eta17-phi7*/	2, 96, 0, 4, 96, 2, 1, 
/* out0158_had-eta18-phi7*/	2, 96, 0, 2, 96, 1, 5, 
/* out0159_had-eta19-phi7*/	1, 96, 1, 2, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 114, 3, 10, 
/* out0162_had-eta2-phi8*/	2, 114, 2, 11, 114, 3, 6, 
/* out0163_had-eta3-phi8*/	2, 113, 3, 13, 114, 2, 5, 
/* out0164_had-eta4-phi8*/	2, 113, 2, 14, 113, 3, 3, 
/* out0165_had-eta5-phi8*/	1, 113, 2, 2, 
/* out0166_had-eta6-phi8*/	2, 52, 0, 5, 70, 2, 10, 
/* out0167_had-eta7-phi8*/	6, 51, 0, 10, 51, 2, 4, 52, 0, 5, 52, 1, 1, 70, 1, 7, 70, 2, 6, 
/* out0168_had-eta8-phi8*/	4, 51, 0, 6, 51, 1, 11, 51, 2, 1, 68, 2, 4, 
/* out0169_had-eta9-phi8*/	3, 49, 0, 1, 68, 1, 4, 68, 2, 12, 
/* out0170_had-eta10-phi8*/	2, 48, 0, 10, 68, 1, 4, 
/* out0171_had-eta11-phi8*/	5, 44, 2, 1, 48, 0, 6, 48, 1, 6, 94, 1, 2, 94, 2, 16, 
/* out0172_had-eta12-phi8*/	4, 44, 2, 10, 48, 1, 1, 94, 1, 5, 99, 0, 6, 
/* out0173_had-eta13-phi8*/	4, 44, 1, 5, 44, 2, 3, 99, 0, 8, 99, 1, 2, 
/* out0174_had-eta14-phi8*/	4, 44, 1, 2, 53, 0, 5, 92, 2, 5, 99, 1, 3, 
/* out0175_had-eta15-phi8*/	4, 53, 0, 5, 53, 1, 1, 92, 1, 1, 92, 2, 6, 
/* out0176_had-eta16-phi8*/	2, 53, 1, 2, 92, 1, 5, 
/* out0177_had-eta17-phi8*/	1, 96, 0, 4, 
/* out0178_had-eta18-phi8*/	1, 96, 0, 4, 
/* out0179_had-eta19-phi8*/	1, 96, 1, 2, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 116, 0, 10, 
/* out0182_had-eta2-phi9*/	2, 116, 0, 6, 116, 1, 11, 
/* out0183_had-eta3-phi9*/	2, 115, 0, 13, 116, 1, 5, 
/* out0184_had-eta4-phi9*/	2, 115, 0, 3, 115, 1, 14, 
/* out0185_had-eta5-phi9*/	1, 115, 1, 2, 
/* out0186_had-eta6-phi9*/	3, 70, 0, 10, 70, 1, 1, 71, 2, 5, 
/* out0187_had-eta7-phi9*/	6, 69, 0, 4, 69, 2, 10, 70, 0, 6, 70, 1, 8, 71, 1, 1, 71, 2, 5, 
/* out0188_had-eta8-phi9*/	4, 68, 0, 4, 69, 0, 1, 69, 1, 11, 69, 2, 6, 
/* out0189_had-eta9-phi9*/	3, 46, 2, 1, 68, 0, 12, 68, 1, 4, 
/* out0190_had-eta10-phi9*/	2, 45, 2, 10, 68, 1, 4, 
/* out0191_had-eta11-phi9*/	5, 44, 0, 1, 45, 1, 6, 45, 2, 6, 94, 0, 16, 94, 1, 3, 
/* out0192_had-eta12-phi9*/	4, 44, 0, 9, 45, 1, 1, 93, 2, 6, 94, 1, 6, 
/* out0193_had-eta13-phi9*/	4, 44, 0, 3, 44, 1, 6, 93, 1, 2, 93, 2, 8, 
/* out0194_had-eta14-phi9*/	4, 39, 2, 5, 44, 1, 2, 92, 0, 5, 93, 1, 3, 
/* out0195_had-eta15-phi9*/	4, 39, 1, 1, 39, 2, 5, 92, 0, 6, 92, 1, 1, 
/* out0196_had-eta16-phi9*/	2, 39, 1, 2, 92, 1, 6, 
/* out0197_had-eta17-phi9*/	2, 92, 1, 1, 105, 2, 4, 
/* out0198_had-eta18-phi9*/	1, 105, 2, 4, 
/* out0199_had-eta19-phi9*/	1, 105, 1, 2, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 116, 3, 10, 
/* out0202_had-eta2-phi10*/	2, 116, 2, 11, 116, 3, 6, 
/* out0203_had-eta3-phi10*/	2, 115, 3, 13, 116, 2, 5, 
/* out0204_had-eta4-phi10*/	2, 115, 2, 14, 115, 3, 3, 
/* out0205_had-eta5-phi10*/	1, 115, 2, 2, 
/* out0206_had-eta6-phi10*/	3, 71, 0, 10, 71, 1, 3, 71, 2, 6, 
/* out0207_had-eta7-phi10*/	3, 47, 2, 7, 69, 0, 7, 71, 1, 12, 
/* out0208_had-eta8-phi10*/	6, 46, 0, 3, 46, 2, 5, 47, 1, 1, 47, 2, 3, 69, 0, 4, 69, 1, 5, 
/* out0209_had-eta9-phi10*/	3, 46, 0, 2, 46, 1, 6, 46, 2, 10, 
/* out0210_had-eta10-phi10*/	3, 45, 0, 11, 46, 1, 4, 95, 2, 2, 
/* out0211_had-eta11-phi10*/	6, 40, 2, 1, 45, 0, 4, 45, 1, 8, 95, 0, 1, 95, 1, 4, 95, 2, 14, 
/* out0212_had-eta12-phi10*/	6, 40, 2, 7, 44, 0, 1, 45, 1, 1, 93, 0, 8, 93, 2, 1, 95, 1, 3, 
/* out0213_had-eta13-phi10*/	9, 39, 0, 1, 39, 2, 1, 40, 1, 2, 40, 2, 3, 44, 0, 2, 44, 1, 1, 93, 0, 4, 93, 1, 5, 93, 2, 1, 
/* out0214_had-eta14-phi10*/	5, 39, 0, 4, 39, 2, 3, 92, 0, 1, 93, 1, 5, 106, 2, 3, 
/* out0215_had-eta15-phi10*/	5, 39, 0, 1, 39, 1, 3, 39, 2, 2, 92, 0, 3, 106, 2, 4, 
/* out0216_had-eta16-phi10*/	7, 39, 1, 5, 92, 0, 1, 92, 1, 1, 105, 0, 2, 105, 2, 2, 106, 1, 1, 106, 2, 1, 
/* out0217_had-eta17-phi10*/	2, 105, 0, 1, 105, 2, 4, 
/* out0218_had-eta18-phi10*/	2, 105, 1, 5, 105, 2, 2, 
/* out0219_had-eta19-phi10*/	1, 105, 1, 2, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 118, 0, 10, 
/* out0222_had-eta2-phi11*/	2, 118, 0, 6, 118, 1, 11, 
/* out0223_had-eta3-phi11*/	2, 117, 0, 13, 118, 1, 5, 
/* out0224_had-eta4-phi11*/	2, 117, 0, 3, 117, 1, 14, 
/* out0225_had-eta5-phi11*/	1, 117, 1, 2, 
/* out0226_had-eta6-phi11*/	1, 71, 0, 5, 
/* out0227_had-eta7-phi11*/	4, 47, 0, 14, 47, 1, 1, 47, 2, 6, 71, 0, 1, 
/* out0228_had-eta8-phi11*/	3, 42, 2, 4, 46, 0, 4, 47, 1, 13, 
/* out0229_had-eta9-phi11*/	5, 41, 0, 1, 41, 2, 1, 42, 2, 4, 46, 0, 7, 46, 1, 5, 
/* out0230_had-eta10-phi11*/	4, 41, 2, 12, 46, 1, 1, 95, 0, 4, 108, 1, 2, 
/* out0231_had-eta11-phi11*/	8, 40, 0, 3, 40, 2, 1, 41, 1, 5, 41, 2, 3, 45, 0, 1, 95, 0, 11, 95, 1, 6, 108, 1, 1, 
/* out0232_had-eta12-phi11*/	6, 40, 0, 6, 40, 1, 1, 40, 2, 4, 93, 0, 1, 95, 1, 3, 107, 2, 8, 
/* out0233_had-eta13-phi11*/	6, 40, 1, 8, 93, 0, 3, 93, 1, 1, 106, 0, 1, 107, 1, 2, 107, 2, 4, 
/* out0234_had-eta14-phi11*/	5, 34, 2, 1, 39, 0, 6, 40, 1, 1, 106, 0, 3, 106, 2, 5, 
/* out0235_had-eta15-phi11*/	4, 39, 0, 4, 39, 1, 2, 106, 1, 3, 106, 2, 3, 
/* out0236_had-eta16-phi11*/	4, 33, 1, 5, 39, 1, 3, 105, 0, 2, 106, 1, 4, 
/* out0237_had-eta17-phi11*/	2, 33, 1, 3, 105, 0, 5, 
/* out0238_had-eta18-phi11*/	2, 105, 0, 2, 105, 1, 5, 
/* out0239_had-eta19-phi11*/	1, 105, 1, 1, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 118, 3, 10, 
/* out0242_had-eta2-phi12*/	2, 118, 2, 11, 118, 3, 6, 
/* out0243_had-eta3-phi12*/	2, 117, 3, 13, 118, 2, 5, 
/* out0244_had-eta4-phi12*/	2, 117, 2, 14, 117, 3, 3, 
/* out0245_had-eta5-phi12*/	1, 117, 2, 2, 
/* out0246_had-eta6-phi12*/	2, 43, 0, 3, 43, 2, 2, 
/* out0247_had-eta7-phi12*/	4, 43, 0, 3, 43, 1, 5, 43, 2, 14, 47, 0, 2, 
/* out0248_had-eta8-phi12*/	4, 42, 0, 11, 42, 2, 6, 43, 1, 3, 47, 1, 1, 
/* out0249_had-eta9-phi12*/	3, 41, 0, 2, 42, 1, 13, 42, 2, 2, 
/* out0250_had-eta10-phi12*/	4, 36, 2, 1, 41, 0, 12, 41, 1, 2, 108, 1, 4, 
/* out0251_had-eta11-phi12*/	6, 35, 2, 3, 40, 0, 1, 41, 1, 9, 107, 0, 2, 108, 0, 8, 108, 1, 9, 
/* out0252_had-eta12-phi12*/	4, 35, 2, 4, 40, 0, 6, 107, 0, 9, 107, 2, 3, 
/* out0253_had-eta13-phi12*/	5, 34, 0, 1, 34, 2, 4, 40, 1, 4, 107, 1, 10, 107, 2, 1, 
/* out0254_had-eta14-phi12*/	4, 34, 2, 7, 90, 2, 1, 106, 0, 8, 107, 1, 1, 
/* out0255_had-eta15-phi12*/	4, 34, 1, 2, 34, 2, 3, 106, 0, 3, 106, 1, 4, 
/* out0256_had-eta16-phi12*/	4, 33, 0, 3, 33, 1, 4, 89, 2, 3, 106, 1, 3, 
/* out0257_had-eta17-phi12*/	4, 33, 0, 1, 33, 1, 4, 89, 2, 3, 105, 0, 2, 
/* out0258_had-eta18-phi12*/	3, 89, 2, 1, 105, 0, 2, 105, 1, 1, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 120, 0, 10, 
/* out0262_had-eta2-phi13*/	2, 120, 0, 6, 120, 1, 11, 
/* out0263_had-eta3-phi13*/	2, 119, 0, 13, 120, 1, 5, 
/* out0264_had-eta4-phi13*/	2, 119, 0, 3, 119, 1, 14, 
/* out0265_had-eta5-phi13*/	1, 119, 1, 2, 
/* out0266_had-eta6-phi13*/	2, 38, 1, 4, 43, 0, 2, 
/* out0267_had-eta7-phi13*/	6, 37, 0, 2, 37, 2, 3, 38, 0, 2, 38, 1, 11, 43, 0, 8, 43, 1, 6, 
/* out0268_had-eta8-phi13*/	5, 37, 0, 1, 37, 1, 2, 37, 2, 13, 42, 0, 4, 43, 1, 2, 
/* out0269_had-eta9-phi13*/	5, 36, 0, 5, 36, 2, 7, 37, 1, 2, 42, 0, 1, 42, 1, 3, 
/* out0270_had-eta10-phi13*/	3, 36, 1, 6, 36, 2, 8, 41, 0, 1, 
/* out0271_had-eta11-phi13*/	4, 35, 0, 7, 35, 2, 5, 91, 2, 6, 108, 0, 8, 
/* out0272_had-eta12-phi13*/	4, 35, 1, 6, 35, 2, 4, 91, 2, 7, 107, 0, 5, 
/* out0273_had-eta13-phi13*/	5, 34, 0, 6, 35, 1, 3, 90, 0, 1, 90, 2, 5, 107, 1, 3, 
/* out0274_had-eta14-phi13*/	4, 34, 0, 3, 34, 1, 2, 34, 2, 1, 90, 2, 8, 
/* out0275_had-eta15-phi13*/	7, 34, 1, 6, 89, 0, 1, 89, 2, 1, 90, 1, 2, 90, 2, 1, 106, 0, 1, 106, 1, 1, 
/* out0276_had-eta16-phi13*/	4, 33, 0, 5, 34, 1, 1, 89, 0, 2, 89, 2, 4, 
/* out0277_had-eta17-phi13*/	3, 33, 0, 3, 89, 1, 1, 89, 2, 4, 
/* out0278_had-eta18-phi13*/	1, 89, 1, 3, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 120, 3, 10, 
/* out0282_had-eta2-phi14*/	2, 120, 2, 11, 120, 3, 6, 
/* out0283_had-eta3-phi14*/	2, 119, 3, 13, 120, 2, 5, 
/* out0284_had-eta4-phi14*/	2, 119, 2, 14, 119, 3, 3, 
/* out0285_had-eta5-phi14*/	1, 119, 2, 2, 
/* out0286_had-eta6-phi14*/	1, 38, 0, 1, 
/* out0287_had-eta7-phi14*/	4, 32, 2, 6, 37, 0, 5, 38, 0, 13, 38, 1, 1, 
/* out0288_had-eta8-phi14*/	4, 31, 2, 2, 32, 2, 1, 37, 0, 8, 37, 1, 10, 
/* out0289_had-eta9-phi14*/	3, 31, 2, 6, 36, 0, 9, 37, 1, 2, 
/* out0290_had-eta10-phi14*/	3, 30, 2, 3, 36, 0, 2, 36, 1, 9, 
/* out0291_had-eta11-phi14*/	5, 30, 2, 5, 35, 0, 7, 36, 1, 1, 91, 0, 11, 91, 2, 1, 
/* out0292_had-eta12-phi14*/	6, 29, 2, 2, 35, 0, 2, 35, 1, 6, 91, 0, 1, 91, 1, 10, 91, 2, 2, 
/* out0293_had-eta13-phi14*/	5, 29, 2, 5, 34, 0, 2, 35, 1, 1, 90, 0, 8, 91, 1, 2, 
/* out0294_had-eta14-phi14*/	6, 29, 2, 1, 34, 0, 4, 34, 1, 2, 90, 0, 3, 90, 1, 5, 90, 2, 1, 
/* out0295_had-eta15-phi14*/	4, 28, 2, 3, 34, 1, 3, 89, 0, 2, 90, 1, 5, 
/* out0296_had-eta16-phi14*/	3, 28, 2, 4, 33, 0, 1, 89, 0, 6, 
/* out0297_had-eta17-phi14*/	4, 28, 2, 1, 33, 0, 3, 89, 0, 1, 89, 1, 4, 
/* out0298_had-eta18-phi14*/	1, 89, 1, 4, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 122, 0, 10, 
/* out0302_had-eta2-phi15*/	2, 122, 0, 6, 122, 1, 11, 
/* out0303_had-eta3-phi15*/	2, 121, 0, 13, 122, 1, 5, 
/* out0304_had-eta4-phi15*/	2, 121, 0, 3, 121, 1, 14, 
/* out0305_had-eta5-phi15*/	1, 121, 1, 2, 
/* out0306_had-eta6-phi15*/	1, 32, 0, 1, 
/* out0307_had-eta7-phi15*/	4, 27, 1, 1, 32, 0, 13, 32, 1, 5, 32, 2, 7, 
/* out0308_had-eta8-phi15*/	4, 31, 0, 10, 31, 2, 2, 32, 1, 8, 32, 2, 2, 
/* out0309_had-eta9-phi15*/	3, 31, 0, 2, 31, 1, 9, 31, 2, 6, 
/* out0310_had-eta10-phi15*/	3, 30, 0, 9, 30, 2, 3, 31, 1, 2, 
/* out0311_had-eta11-phi15*/	6, 30, 0, 1, 30, 1, 7, 30, 2, 5, 88, 0, 2, 88, 1, 16, 91, 0, 3, 
/* out0312_had-eta12-phi15*/	7, 29, 0, 6, 29, 2, 2, 30, 1, 2, 87, 0, 2, 87, 2, 6, 91, 0, 1, 91, 1, 4, 
/* out0313_had-eta13-phi15*/	5, 29, 0, 1, 29, 1, 3, 29, 2, 5, 87, 2, 8, 90, 0, 2, 
/* out0314_had-eta14-phi15*/	9, 28, 0, 2, 29, 1, 4, 29, 2, 1, 86, 0, 1, 86, 2, 2, 87, 1, 1, 87, 2, 1, 90, 0, 2, 90, 1, 3, 
/* out0315_had-eta15-phi15*/	4, 28, 0, 3, 28, 2, 3, 86, 2, 6, 90, 1, 1, 
/* out0316_had-eta16-phi15*/	4, 28, 1, 1, 28, 2, 4, 86, 2, 3, 89, 0, 3, 
/* out0317_had-eta17-phi15*/	5, 28, 1, 3, 28, 2, 1, 85, 1, 2, 89, 0, 1, 89, 1, 3, 
/* out0318_had-eta18-phi15*/	2, 85, 1, 6, 89, 1, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 122, 3, 10, 
/* out0322_had-eta2-phi16*/	2, 122, 2, 11, 122, 3, 6, 
/* out0323_had-eta3-phi16*/	2, 121, 3, 13, 122, 2, 5, 
/* out0324_had-eta4-phi16*/	2, 121, 2, 14, 121, 3, 3, 
/* out0325_had-eta5-phi16*/	1, 121, 2, 2, 
/* out0326_had-eta6-phi16*/	2, 27, 0, 2, 27, 1, 4, 
/* out0327_had-eta7-phi16*/	6, 26, 0, 6, 26, 2, 3, 27, 0, 8, 27, 1, 11, 32, 0, 2, 32, 1, 2, 
/* out0328_had-eta8-phi16*/	5, 26, 0, 2, 26, 1, 4, 26, 2, 13, 31, 0, 2, 32, 1, 1, 
/* out0329_had-eta9-phi16*/	5, 25, 0, 3, 25, 2, 7, 26, 1, 1, 31, 0, 2, 31, 1, 5, 
/* out0330_had-eta10-phi16*/	3, 25, 1, 1, 25, 2, 8, 30, 0, 6, 
/* out0331_had-eta11-phi16*/	4, 24, 2, 5, 30, 1, 7, 84, 2, 1, 88, 0, 13, 
/* out0332_had-eta12-phi16*/	3, 24, 2, 4, 29, 0, 6, 87, 0, 11, 
/* out0333_had-eta13-phi16*/	4, 29, 0, 3, 29, 1, 6, 87, 1, 8, 87, 2, 1, 
/* out0334_had-eta14-phi16*/	5, 23, 2, 1, 28, 0, 2, 29, 1, 3, 86, 0, 6, 87, 1, 2, 
/* out0335_had-eta15-phi16*/	4, 28, 0, 6, 86, 0, 2, 86, 1, 1, 86, 2, 3, 
/* out0336_had-eta16-phi16*/	4, 28, 0, 1, 28, 1, 5, 86, 1, 5, 86, 2, 2, 
/* out0337_had-eta17-phi16*/	3, 28, 1, 3, 85, 0, 4, 85, 1, 2, 
/* out0338_had-eta18-phi16*/	1, 85, 1, 6, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 124, 0, 10, 
/* out0342_had-eta2-phi17*/	2, 124, 0, 6, 124, 1, 11, 
/* out0343_had-eta3-phi17*/	2, 123, 0, 13, 124, 1, 5, 
/* out0344_had-eta4-phi17*/	2, 123, 0, 3, 123, 1, 14, 
/* out0345_had-eta5-phi17*/	1, 123, 1, 2, 
/* out0346_had-eta6-phi17*/	3, 21, 0, 4, 21, 2, 2, 27, 0, 3, 
/* out0347_had-eta7-phi17*/	5, 21, 0, 2, 21, 1, 2, 21, 2, 14, 26, 0, 5, 27, 0, 3, 
/* out0348_had-eta8-phi17*/	4, 19, 0, 1, 19, 2, 6, 26, 0, 3, 26, 1, 11, 
/* out0349_had-eta9-phi17*/	3, 19, 2, 2, 25, 0, 13, 25, 1, 2, 
/* out0350_had-eta10-phi17*/	4, 24, 0, 2, 25, 1, 12, 25, 2, 1, 84, 0, 2, 
/* out0351_had-eta11-phi17*/	6, 24, 0, 9, 24, 1, 1, 24, 2, 3, 84, 0, 5, 84, 2, 9, 88, 0, 1, 
/* out0352_had-eta12-phi17*/	7, 24, 1, 6, 24, 2, 4, 82, 0, 1, 84, 1, 3, 84, 2, 6, 87, 0, 3, 87, 1, 1, 
/* out0353_had-eta13-phi17*/	4, 23, 0, 4, 23, 2, 4, 82, 2, 6, 87, 1, 4, 
/* out0354_had-eta14-phi17*/	3, 23, 2, 7, 82, 2, 4, 86, 0, 4, 
/* out0355_had-eta15-phi17*/	4, 23, 2, 3, 28, 0, 2, 86, 0, 3, 86, 1, 4, 
/* out0356_had-eta16-phi17*/	4, 22, 2, 3, 28, 1, 3, 81, 2, 1, 86, 1, 5, 
/* out0357_had-eta17-phi17*/	3, 22, 2, 3, 28, 1, 1, 85, 0, 5, 
/* out0358_had-eta18-phi17*/	1, 85, 0, 3, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 124, 3, 10, 
/* out0362_had-eta2-phi18*/	2, 124, 2, 11, 124, 3, 6, 
/* out0363_had-eta3-phi18*/	2, 123, 3, 13, 124, 2, 5, 
/* out0364_had-eta4-phi18*/	2, 123, 2, 14, 123, 3, 3, 
/* out0365_had-eta5-phi18*/	1, 123, 2, 2, 
/* out0366_had-eta6-phi18*/	1, 21, 0, 2, 
/* out0367_had-eta7-phi18*/	4, 19, 0, 1, 20, 2, 6, 21, 0, 8, 21, 1, 14, 
/* out0368_had-eta8-phi18*/	3, 19, 0, 13, 19, 1, 4, 19, 2, 4, 
/* out0369_had-eta9-phi18*/	5, 17, 0, 5, 17, 2, 1, 19, 1, 7, 19, 2, 4, 25, 1, 1, 
/* out0370_had-eta10-phi18*/	3, 17, 0, 1, 17, 2, 12, 84, 0, 2, 
/* out0371_had-eta11-phi18*/	7, 16, 2, 1, 17, 1, 1, 17, 2, 3, 24, 0, 5, 24, 1, 3, 84, 0, 7, 84, 1, 6, 
/* out0372_had-eta12-phi18*/	6, 16, 2, 4, 23, 0, 1, 24, 1, 6, 82, 0, 4, 83, 2, 1, 84, 1, 7, 
/* out0373_had-eta13-phi18*/	4, 23, 0, 8, 82, 0, 7, 82, 1, 1, 82, 2, 3, 
/* out0374_had-eta14-phi18*/	5, 23, 0, 1, 23, 1, 6, 23, 2, 1, 82, 1, 5, 82, 2, 3, 
/* out0375_had-eta15-phi18*/	6, 22, 0, 2, 23, 1, 4, 81, 0, 3, 81, 2, 3, 82, 1, 1, 86, 1, 1, 
/* out0376_had-eta16-phi18*/	3, 22, 0, 3, 22, 2, 3, 81, 2, 6, 
/* out0377_had-eta17-phi18*/	3, 22, 2, 6, 81, 2, 3, 85, 0, 2, 
/* out0378_had-eta18-phi18*/	1, 85, 0, 2, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 126, 0, 10, 
/* out0382_had-eta2-phi19*/	2, 126, 0, 6, 126, 1, 11, 
/* out0383_had-eta3-phi19*/	2, 125, 0, 13, 126, 1, 5, 
/* out0384_had-eta4-phi19*/	2, 125, 0, 3, 125, 1, 14, 
/* out0385_had-eta5-phi19*/	1, 125, 1, 2, 
/* out0386_had-eta6-phi19*/	1, 20, 0, 3, 
/* out0387_had-eta7-phi19*/	3, 20, 0, 12, 20, 1, 7, 20, 2, 7, 
/* out0388_had-eta8-phi19*/	6, 18, 0, 5, 18, 2, 5, 19, 0, 1, 19, 1, 3, 20, 1, 4, 20, 2, 3, 
/* out0389_had-eta9-phi19*/	3, 17, 0, 6, 18, 2, 10, 19, 1, 2, 
/* out0390_had-eta10-phi19*/	2, 17, 0, 4, 17, 1, 11, 
/* out0391_had-eta11-phi19*/	5, 16, 0, 8, 16, 2, 1, 17, 1, 4, 83, 0, 8, 83, 2, 4, 
/* out0392_had-eta12-phi19*/	6, 16, 0, 1, 16, 1, 1, 16, 2, 7, 82, 0, 1, 83, 1, 1, 83, 2, 10, 
/* out0393_had-eta13-phi19*/	10, 11, 2, 1, 16, 1, 2, 16, 2, 3, 23, 0, 2, 23, 1, 1, 79, 2, 1, 82, 0, 3, 82, 1, 4, 83, 1, 1, 83, 2, 1, 
/* out0394_had-eta14-phi19*/	5, 11, 2, 3, 23, 1, 4, 79, 2, 2, 81, 0, 1, 82, 1, 5, 
/* out0395_had-eta15-phi19*/	4, 11, 2, 1, 22, 0, 3, 23, 1, 1, 81, 0, 7, 
/* out0396_had-eta16-phi19*/	4, 22, 0, 5, 81, 0, 1, 81, 1, 3, 81, 2, 2, 
/* out0397_had-eta17-phi19*/	4, 22, 1, 5, 22, 2, 1, 81, 1, 3, 81, 2, 1, 
/* out0398_had-eta18-phi19*/	1, 22, 1, 1, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 126, 3, 10, 
/* out0402_had-eta2-phi20*/	2, 126, 2, 11, 126, 3, 6, 
/* out0403_had-eta3-phi20*/	2, 125, 3, 13, 126, 2, 5, 
/* out0404_had-eta4-phi20*/	2, 125, 2, 14, 125, 3, 3, 
/* out0405_had-eta5-phi20*/	1, 125, 2, 2, 
/* out0406_had-eta6-phi20*/	0, 
/* out0407_had-eta7-phi20*/	4, 20, 0, 1, 20, 1, 4, 67, 0, 7, 67, 2, 10, 
/* out0408_had-eta8-phi20*/	4, 18, 0, 11, 18, 1, 4, 20, 1, 1, 67, 2, 6, 
/* out0409_had-eta9-phi20*/	3, 18, 1, 12, 18, 2, 1, 64, 0, 4, 
/* out0410_had-eta10-phi20*/	2, 64, 0, 4, 64, 2, 10, 
/* out0411_had-eta11-phi20*/	5, 16, 0, 6, 16, 1, 1, 64, 2, 6, 83, 0, 8, 83, 1, 2, 
/* out0412_had-eta12-phi20*/	4, 16, 0, 1, 16, 1, 9, 79, 0, 1, 83, 1, 11, 
/* out0413_had-eta13-phi20*/	5, 11, 0, 5, 16, 1, 3, 79, 0, 7, 79, 2, 3, 83, 1, 1, 
/* out0414_had-eta14-phi20*/	3, 11, 0, 2, 11, 2, 5, 79, 2, 8, 
/* out0415_had-eta15-phi20*/	5, 11, 2, 6, 22, 0, 1, 79, 2, 2, 81, 0, 4, 81, 1, 1, 
/* out0416_had-eta16-phi20*/	3, 22, 0, 2, 22, 1, 3, 81, 1, 6, 
/* out0417_had-eta17-phi20*/	2, 22, 1, 5, 81, 1, 3, 
/* out0418_had-eta18-phi20*/	1, 22, 1, 2, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 128, 0, 10, 
/* out0422_had-eta2-phi21*/	2, 128, 0, 6, 128, 1, 11, 
/* out0423_had-eta3-phi21*/	2, 127, 0, 13, 128, 1, 5, 
/* out0424_had-eta4-phi21*/	2, 127, 0, 3, 127, 1, 14, 
/* out0425_had-eta5-phi21*/	1, 127, 1, 2, 
/* out0426_had-eta6-phi21*/	1, 67, 0, 1, 
/* out0427_had-eta7-phi21*/	4, 66, 0, 1, 66, 2, 4, 67, 0, 8, 67, 1, 10, 
/* out0428_had-eta8-phi21*/	4, 65, 0, 11, 65, 2, 4, 66, 2, 1, 67, 1, 6, 
/* out0429_had-eta9-phi21*/	3, 64, 0, 4, 65, 1, 1, 65, 2, 12, 
/* out0430_had-eta10-phi21*/	2, 64, 0, 4, 64, 1, 10, 
/* out0431_had-eta11-phi21*/	5, 12, 0, 6, 12, 2, 1, 64, 1, 6, 80, 0, 8, 80, 2, 2, 
/* out0432_had-eta12-phi21*/	4, 12, 0, 1, 12, 2, 9, 79, 0, 1, 80, 2, 11, 
/* out0433_had-eta13-phi21*/	5, 11, 0, 6, 12, 2, 3, 79, 0, 7, 79, 1, 2, 80, 2, 1, 
/* out0434_had-eta14-phi21*/	3, 11, 0, 2, 11, 1, 5, 79, 1, 8, 
/* out0435_had-eta15-phi21*/	5, 5, 0, 1, 11, 1, 5, 76, 0, 4, 76, 2, 1, 79, 1, 2, 
/* out0436_had-eta16-phi21*/	3, 5, 0, 2, 5, 2, 3, 76, 2, 6, 
/* out0437_had-eta17-phi21*/	2, 5, 2, 5, 76, 2, 3, 
/* out0438_had-eta18-phi21*/	1, 5, 2, 2, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 128, 3, 10, 
/* out0442_had-eta2-phi22*/	2, 128, 2, 11, 128, 3, 6, 
/* out0443_had-eta3-phi22*/	2, 127, 3, 13, 128, 2, 5, 
/* out0444_had-eta4-phi22*/	2, 127, 2, 14, 127, 3, 3, 
/* out0445_had-eta5-phi22*/	1, 127, 2, 2, 
/* out0446_had-eta6-phi22*/	1, 66, 0, 3, 
/* out0447_had-eta7-phi22*/	3, 66, 0, 12, 66, 1, 7, 66, 2, 7, 
/* out0448_had-eta8-phi22*/	6, 14, 0, 1, 14, 2, 3, 65, 0, 5, 65, 1, 5, 66, 1, 3, 66, 2, 4, 
/* out0449_had-eta9-phi22*/	3, 13, 0, 6, 14, 2, 2, 65, 1, 10, 
/* out0450_had-eta10-phi22*/	2, 13, 0, 4, 13, 2, 11, 
/* out0451_had-eta11-phi22*/	5, 12, 0, 8, 12, 1, 1, 13, 2, 4, 80, 0, 8, 80, 1, 4, 
/* out0452_had-eta12-phi22*/	6, 12, 0, 1, 12, 1, 7, 12, 2, 1, 77, 0, 1, 80, 1, 10, 80, 2, 1, 
/* out0453_had-eta13-phi22*/	11, 6, 0, 2, 6, 2, 1, 11, 0, 1, 11, 1, 1, 12, 1, 3, 12, 2, 2, 77, 0, 3, 77, 2, 4, 79, 1, 2, 80, 1, 1, 80, 2, 1, 
/* out0454_had-eta14-phi22*/	5, 6, 2, 4, 11, 1, 3, 76, 0, 1, 77, 2, 5, 79, 1, 2, 
/* out0455_had-eta15-phi22*/	4, 5, 0, 3, 6, 2, 1, 11, 1, 2, 76, 0, 7, 
/* out0456_had-eta16-phi22*/	4, 5, 0, 5, 76, 0, 1, 76, 1, 2, 76, 2, 3, 
/* out0457_had-eta17-phi22*/	4, 5, 1, 1, 5, 2, 5, 76, 1, 1, 76, 2, 3, 
/* out0458_had-eta18-phi22*/	1, 5, 2, 1, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 130, 0, 10, 
/* out0462_had-eta2-phi23*/	2, 130, 0, 6, 130, 1, 11, 
/* out0463_had-eta3-phi23*/	2, 129, 0, 13, 130, 1, 5, 
/* out0464_had-eta4-phi23*/	2, 129, 0, 3, 129, 1, 14, 
/* out0465_had-eta5-phi23*/	1, 129, 1, 2, 
/* out0466_had-eta6-phi23*/	1, 15, 0, 2, 
/* out0467_had-eta7-phi23*/	4, 14, 0, 1, 15, 0, 8, 15, 2, 14, 66, 1, 6, 
/* out0468_had-eta8-phi23*/	3, 14, 0, 13, 14, 1, 4, 14, 2, 4, 
/* out0469_had-eta9-phi23*/	5, 8, 2, 1, 13, 0, 5, 13, 1, 1, 14, 1, 4, 14, 2, 7, 
/* out0470_had-eta10-phi23*/	3, 13, 0, 1, 13, 1, 12, 78, 0, 2, 
/* out0471_had-eta11-phi23*/	7, 7, 0, 5, 7, 2, 3, 12, 1, 1, 13, 1, 3, 13, 2, 1, 78, 0, 7, 78, 2, 6, 
/* out0472_had-eta12-phi23*/	6, 6, 0, 1, 7, 2, 6, 12, 1, 4, 77, 0, 4, 78, 2, 7, 80, 1, 1, 
/* out0473_had-eta13-phi23*/	4, 6, 0, 8, 77, 0, 7, 77, 1, 3, 77, 2, 1, 
/* out0474_had-eta14-phi23*/	5, 6, 0, 1, 6, 1, 1, 6, 2, 6, 77, 1, 3, 77, 2, 5, 
/* out0475_had-eta15-phi23*/	6, 5, 0, 2, 6, 2, 4, 73, 2, 1, 76, 0, 3, 76, 1, 3, 77, 2, 1, 
/* out0476_had-eta16-phi23*/	3, 5, 0, 3, 5, 1, 3, 76, 1, 6, 
/* out0477_had-eta17-phi23*/	3, 5, 1, 6, 72, 0, 2, 76, 1, 3, 
/* out0478_had-eta18-phi23*/	1, 72, 0, 2, 
/* out0479_had-eta19-phi23*/	0, 
};