parameter integer matrixH [0:7328] = {
/* num inputs = 140(in0-in139) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 13 */
//* total number of input in adders 2282 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	6,114,1,16,114,2,8,115,0,3,115,1,2,125,1,2,125,2,12,
/* out0004_em-eta4-phi0*/	6,102,1,16,102,2,6,103,1,1,114,2,8,115,0,12,115,2,1,
/* out0005_em-eta5-phi0*/	3,90,1,9,102,2,10,103,0,10,
/* out0006_em-eta6-phi0*/	4,90,1,7,90,2,14,91,0,3,103,0,1,
/* out0007_em-eta7-phi0*/	3,78,1,12,90,2,2,91,0,4,
/* out0008_em-eta8-phi0*/	5,78,1,1,78,2,12,79,0,2,214,0,9,214,1,1,
/* out0009_em-eta9-phi0*/	6,62,1,11,78,2,3,79,0,1,214,0,7,214,1,6,214,2,6,
/* out0010_em-eta10-phi0*/	6,62,1,1,62,2,12,63,0,1,205,0,8,205,1,1,214,2,7,
/* out0011_em-eta11-phi0*/	9,44,4,15,44,5,2,45,0,5,45,1,16,62,2,2,63,0,3,205,0,4,205,1,3,205,2,6,
/* out0012_em-eta12-phi0*/	6,44,5,6,45,0,11,45,4,8,45,5,3,196,0,6,205,2,6,
/* out0013_em-eta13-phi0*/	7,45,2,12,45,3,4,45,4,8,45,5,4,196,0,6,196,1,1,196,2,3,
/* out0014_em-eta14-phi0*/	8,26,4,12,26,5,1,27,0,1,27,1,16,45,2,2,45,3,12,187,0,1,196,2,8,
/* out0015_em-eta15-phi0*/	5,26,5,3,27,0,12,27,4,3,187,0,7,196,2,2,
/* out0016_em-eta16-phi0*/	6,27,2,1,27,3,13,27,4,10,27,5,2,187,0,3,187,2,3,
/* out0017_em-eta17-phi0*/	4,12,3,2,27,2,8,27,3,3,187,2,5,
/* out0018_em-eta18-phi0*/	5,11,2,10,11,3,4,12,3,12,12,4,4,187,2,2,
/* out0019_em-eta19-phi0*/	5,11,0,5,11,1,16,11,2,6,11,3,1,12,4,12,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	1,126,1,1,
/* out0023_em-eta3-phi1*/	5,115,1,9,125,1,14,125,2,4,126,0,14,126,1,1,
/* out0024_em-eta4-phi1*/	5,103,1,3,115,0,1,115,1,5,115,2,15,116,0,6,
/* out0025_em-eta5-phi1*/	4,103,0,4,103,1,11,103,2,10,116,0,1,
/* out0026_em-eta6-phi1*/	5,91,0,3,91,1,12,103,0,1,103,2,5,104,0,1,
/* out0027_em-eta7-phi1*/	5,78,1,1,79,1,1,91,0,6,91,1,1,91,2,11,
/* out0028_em-eta8-phi1*/	7,78,1,2,78,2,1,79,0,7,79,1,7,214,1,1,222,1,1,222,2,9,
/* out0029_em-eta9-phi1*/	8,62,1,1,64,1,1,79,0,6,79,2,5,214,1,7,215,0,6,222,1,3,222,2,4,
/* out0030_em-eta10-phi1*/	13,62,1,3,62,2,2,63,0,3,63,1,15,63,2,5,64,0,2,64,1,11,205,0,4,205,1,3,214,1,1,214,2,3,215,0,4,215,2,7,
/* out0031_em-eta11-phi1*/	11,44,4,1,44,5,1,63,0,9,63,1,1,63,2,9,63,3,12,64,3,1,205,1,8,205,2,3,206,0,3,215,2,1,
/* out0032_em-eta12-phi1*/	12,44,5,7,45,5,7,46,1,4,47,1,2,63,3,4,64,3,3,196,0,2,196,1,2,205,1,1,205,2,1,206,0,2,206,2,3,
/* out0033_em-eta13-phi1*/	7,45,2,2,45,5,2,46,0,8,46,1,10,46,2,1,196,0,2,196,1,9,
/* out0034_em-eta14-phi1*/	8,26,4,4,26,5,1,46,0,8,46,3,6,187,0,1,196,1,3,196,2,3,197,0,1,
/* out0035_em-eta15-phi1*/	7,26,5,11,27,0,3,27,4,1,27,5,4,46,3,1,187,0,3,187,1,4,
/* out0036_em-eta16-phi1*/	8,27,2,2,27,4,2,27,5,9,28,0,1,28,1,1,187,0,1,187,1,5,187,2,1,
/* out0037_em-eta17-phi1*/	5,12,3,1,27,2,5,28,0,6,187,1,1,187,2,3,
/* out0038_em-eta18-phi1*/	5,11,0,2,11,3,11,12,3,1,28,0,2,187,2,1,
/* out0039_em-eta19-phi1*/	1,11,0,6,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	4,126,1,2,134,0,4,134,1,1,134,2,2,
/* out0043_em-eta3-phi2*/	7,126,0,2,126,1,12,126,2,15,127,0,5,134,0,9,134,1,9,134,2,5,
/* out0044_em-eta4-phi2*/	5,116,0,7,116,1,15,116,2,7,126,2,1,127,0,2,
/* out0045_em-eta5-phi2*/	6,103,1,1,103,2,1,104,0,5,104,1,10,116,0,2,116,2,7,
/* out0046_em-eta6-phi2*/	4,91,1,3,92,1,1,104,0,10,104,2,6,
/* out0047_em-eta7-phi2*/	4,79,1,1,91,2,5,92,0,10,92,1,2,
/* out0048_em-eta8-phi2*/	7,79,1,7,79,2,3,80,0,1,92,0,4,222,1,7,222,2,3,223,0,8,
/* out0049_em-eta9-phi2*/	8,63,4,5,79,2,8,80,0,3,215,0,5,215,1,6,222,1,5,223,0,4,223,2,3,
/* out0050_em-eta10-phi2*/	9,63,4,11,63,5,9,64,0,14,64,1,4,64,4,1,64,5,1,215,0,1,215,1,8,215,2,6,
/* out0051_em-eta11-phi2*/	8,63,2,2,64,2,5,64,3,6,64,4,15,64,5,4,206,0,9,206,1,2,215,2,2,
/* out0052_em-eta12-phi2*/	7,46,4,6,47,1,13,64,2,4,64,3,6,206,0,2,206,1,2,206,2,7,
/* out0053_em-eta13-phi2*/	8,46,1,2,46,2,10,47,0,10,47,1,1,47,4,1,196,1,1,197,0,5,206,2,4,
/* out0054_em-eta14-phi2*/	6,46,2,5,46,3,6,47,3,4,47,4,5,197,0,6,197,2,2,
/* out0055_em-eta15-phi2*/	7,27,5,1,28,1,1,29,1,5,46,3,3,47,3,6,187,1,1,197,2,5,
/* out0056_em-eta16-phi2*/	5,28,1,11,28,2,1,29,1,2,187,1,3,188,1,1,
/* out0057_em-eta17-phi2*/	6,28,0,4,28,1,3,28,2,3,28,3,1,187,1,2,188,1,2,
/* out0058_em-eta18-phi2*/	4,28,0,3,28,3,6,187,2,1,188,1,1,
/* out0059_em-eta19-phi2*/	2,11,0,3,28,3,3,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	7,127,0,5,127,1,16,127,2,7,134,0,3,134,1,6,134,2,9,135,2,6,
/* out0064_em-eta4-phi3*/	6,116,1,1,116,2,2,117,0,6,117,1,10,127,0,4,127,2,8,
/* out0065_em-eta5-phi3*/	6,104,1,6,104,2,2,105,0,1,105,1,2,117,0,10,117,2,5,
/* out0066_em-eta6-phi3*/	3,92,1,4,104,2,8,105,0,9,
/* out0067_em-eta7-phi3*/	3,92,0,2,92,1,9,92,2,7,
/* out0068_em-eta8-phi3*/	5,80,0,1,80,1,6,92,2,7,223,0,2,223,1,7,
/* out0069_em-eta9-phi3*/	7,80,0,8,80,1,2,80,2,2,216,0,2,223,0,2,223,1,4,223,2,12,
/* out0070_em-eta10-phi3*/	9,63,5,7,64,5,4,65,1,2,66,1,4,80,0,3,80,2,2,215,1,2,216,0,12,216,2,2,
/* out0071_em-eta11-phi3*/	6,64,2,6,64,5,7,65,0,8,65,1,13,206,1,5,216,2,7,
/* out0072_em-eta12-phi3*/	8,46,4,10,46,5,5,64,2,1,65,0,8,65,3,3,206,1,7,206,2,1,207,0,3,
/* out0073_em-eta13-phi3*/	8,46,5,7,47,0,6,47,4,5,47,5,5,197,0,3,197,1,3,206,2,1,207,2,1,
/* out0074_em-eta14-phi3*/	7,47,2,8,47,3,4,47,4,5,47,5,3,197,0,1,197,1,5,197,2,2,
/* out0075_em-eta15-phi3*/	5,28,4,6,29,1,5,47,2,3,47,3,2,197,2,6,
/* out0076_em-eta16-phi3*/	5,28,2,2,29,0,8,29,1,4,188,1,1,188,2,4,
/* out0077_em-eta17-phi3*/	4,28,2,8,29,0,1,29,4,2,188,1,4,
/* out0078_em-eta18-phi3*/	5,28,2,2,28,3,3,29,3,2,29,4,2,188,1,2,
/* out0079_em-eta19-phi3*/	2,28,3,3,29,3,5,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	3,135,1,3,135,2,4,136,0,3,
/* out0083_em-eta3-phi4*/	8,127,2,1,128,0,5,128,1,13,128,2,1,135,1,13,135,2,6,136,0,3,136,2,1,
/* out0084_em-eta4-phi4*/	6,117,1,6,117,2,3,118,0,2,118,1,3,128,0,11,128,2,7,
/* out0085_em-eta5-phi4*/	3,105,1,9,117,2,8,118,0,9,
/* out0086_em-eta6-phi4*/	3,105,0,5,105,1,5,105,2,11,
/* out0087_em-eta7-phi4*/	5,92,2,2,93,0,6,93,1,6,105,0,1,105,2,2,
/* out0088_em-eta8-phi4*/	5,80,1,5,93,0,10,223,1,2,224,0,2,224,1,2,
/* out0089_em-eta9-phi4*/	10,80,1,3,80,2,8,81,0,1,216,0,1,216,1,1,223,1,3,223,2,1,224,0,14,224,1,1,224,2,6,
/* out0090_em-eta10-phi4*/	9,65,4,12,65,5,1,66,0,1,66,1,10,80,2,4,216,0,1,216,1,13,216,2,1,224,2,1,
/* out0091_em-eta11-phi4*/	9,65,1,1,65,2,13,66,0,13,66,1,2,66,4,5,207,0,5,207,1,1,216,1,2,216,2,6,
/* out0092_em-eta12-phi4*/	8,46,5,1,65,2,3,65,3,12,66,3,9,66,4,3,207,0,8,207,1,1,207,2,2,
/* out0093_em-eta13-phi4*/	8,46,5,3,47,5,7,48,1,8,49,1,4,65,3,1,66,3,1,197,1,1,207,2,8,
/* out0094_em-eta14-phi4*/	6,47,2,5,47,5,1,48,0,9,48,1,4,197,1,5,198,0,3,
/* out0095_em-eta15-phi4*/	8,28,4,10,28,5,1,48,0,5,188,2,2,197,1,2,197,2,1,198,0,2,198,2,1,
/* out0096_em-eta16-phi4*/	3,28,5,7,29,0,6,188,2,6,
/* out0097_em-eta17-phi4*/	6,29,0,1,29,4,10,29,5,1,188,0,2,188,1,2,188,2,1,
/* out0098_em-eta18-phi4*/	4,29,2,2,29,3,5,29,4,2,188,1,2,
/* out0099_em-eta19-phi4*/	2,29,2,1,29,3,4,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	1,136,0,2,
/* out0103_em-eta3-phi5*/	6,128,1,3,128,2,3,129,0,3,129,1,8,136,0,8,136,2,15,
/* out0104_em-eta4-phi5*/	4,118,1,12,118,2,1,128,2,5,129,0,13,
/* out0105_em-eta5-phi5*/	4,106,1,4,118,0,5,118,1,1,118,2,15,
/* out0106_em-eta6-phi5*/	3,105,2,3,106,0,13,106,1,4,
/* out0107_em-eta7-phi5*/	3,93,1,10,93,2,5,106,0,3,
/* out0108_em-eta8-phi5*/	3,81,1,4,93,2,11,224,1,3,
/* out0109_em-eta9-phi5*/	5,81,0,8,81,1,4,217,0,1,224,1,10,224,2,7,
/* out0110_em-eta10-phi5*/	5,65,4,4,65,5,9,81,0,7,217,0,13,224,2,2,
/* out0111_em-eta11-phi5*/	8,65,5,6,66,0,2,66,2,3,66,4,7,66,5,16,207,1,3,217,0,2,217,2,8,
/* out0112_em-eta12-phi5*/	6,48,4,6,49,1,1,66,2,13,66,3,6,66,4,1,207,1,10,
/* out0113_em-eta13-phi5*/	8,48,1,2,48,2,1,48,4,2,49,0,7,49,1,11,198,0,3,207,1,1,207,2,5,
/* out0114_em-eta14-phi5*/	6,48,0,1,48,1,2,48,2,14,48,3,2,49,0,1,198,0,7,
/* out0115_em-eta15-phi5*/	6,28,5,1,48,0,1,48,2,1,48,3,13,198,0,1,198,2,5,
/* out0116_em-eta16-phi5*/	6,28,5,7,29,5,6,48,3,1,188,0,1,188,2,3,198,2,2,
/* out0117_em-eta17-phi5*/	3,29,2,3,29,5,9,188,0,10,
/* out0118_em-eta18-phi5*/	3,29,2,9,188,0,3,188,1,1,
/* out0119_em-eta19-phi5*/	1,29,2,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	1,137,2,2,
/* out0123_em-eta3-phi6*/	6,129,1,8,129,2,3,130,0,3,130,1,3,137,1,9,137,2,14,
/* out0124_em-eta4-phi6*/	4,119,0,1,119,1,12,129,2,13,130,0,5,
/* out0125_em-eta5-phi6*/	4,106,1,4,119,0,15,119,1,1,119,2,5,
/* out0126_em-eta6-phi6*/	3,106,1,4,106,2,13,107,0,3,
/* out0127_em-eta7-phi6*/	3,94,0,5,94,1,10,106,2,3,
/* out0128_em-eta8-phi6*/	4,81,1,4,94,0,11,225,0,1,225,1,3,
/* out0129_em-eta9-phi6*/	6,81,1,4,81,2,8,217,1,1,225,0,15,225,1,3,225,2,8,
/* out0130_em-eta10-phi6*/	5,67,4,4,68,1,9,81,2,7,217,1,13,225,2,2,
/* out0131_em-eta11-phi6*/	8,67,0,3,67,1,16,67,2,7,68,0,2,68,1,6,208,0,3,217,1,2,217,2,8,
/* out0132_em-eta12-phi6*/	6,48,4,6,48,5,1,67,0,13,67,2,1,67,3,6,208,0,10,
/* out0133_em-eta13-phi6*/	8,48,4,2,48,5,11,49,0,7,49,4,1,49,5,2,198,1,3,208,0,1,208,2,5,
/* out0134_em-eta14-phi6*/	6,49,0,1,49,2,1,49,3,2,49,4,14,49,5,2,198,1,7,
/* out0135_em-eta15-phi6*/	6,31,1,1,49,2,1,49,3,13,49,4,1,198,1,1,198,2,5,
/* out0136_em-eta16-phi6*/	6,30,1,6,31,1,7,49,3,1,189,1,1,189,2,3,198,2,2,
/* out0137_em-eta17-phi6*/	3,30,0,3,30,1,9,189,1,4,
/* out0138_em-eta18-phi6*/	2,30,0,9,189,1,2,
/* out0139_em-eta19-phi6*/	1,30,0,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	2,137,1,2,138,0,7,
/* out0143_em-eta3-phi7*/	7,130,0,1,130,1,13,130,2,5,131,0,1,137,1,5,138,0,8,138,2,12,
/* out0144_em-eta4-phi7*/	6,119,1,3,119,2,2,120,0,3,120,1,6,130,0,7,130,2,11,
/* out0145_em-eta5-phi7*/	3,107,1,9,119,2,9,120,0,8,
/* out0146_em-eta6-phi7*/	3,107,0,11,107,1,5,107,2,5,
/* out0147_em-eta7-phi7*/	5,94,1,6,94,2,6,95,0,2,107,0,2,107,2,1,
/* out0148_em-eta8-phi7*/	5,82,1,5,94,2,10,225,1,3,226,0,3,226,1,1,
/* out0149_em-eta9-phi7*/	8,81,2,1,82,0,8,82,1,3,218,0,1,218,1,1,225,1,7,225,2,5,226,0,7,
/* out0150_em-eta10-phi7*/	9,67,4,12,67,5,10,68,0,1,68,1,1,82,0,4,218,0,13,218,1,1,218,2,1,225,2,1,
/* out0151_em-eta11-phi7*/	9,67,2,5,67,5,2,68,0,13,68,4,13,68,5,1,208,0,1,208,1,5,218,0,2,218,2,6,
/* out0152_em-eta12-phi7*/	8,51,1,1,67,2,3,67,3,9,68,3,12,68,4,3,208,0,1,208,1,8,208,2,2,
/* out0153_em-eta13-phi7*/	8,48,5,4,49,5,8,50,1,7,51,1,3,67,3,1,68,3,1,199,0,1,208,2,8,
/* out0154_em-eta14-phi7*/	6,49,2,9,49,5,4,50,0,5,50,1,1,198,1,3,199,0,5,
/* out0155_em-eta15-phi7*/	8,30,4,10,31,1,1,49,2,5,189,2,1,198,1,2,198,2,1,199,0,2,199,2,1,
/* out0156_em-eta16-phi7*/	3,31,0,6,31,1,7,189,2,6,
/* out0157_em-eta17-phi7*/	5,30,1,1,30,2,10,31,0,1,189,1,3,189,2,1,
/* out0158_em-eta18-phi7*/	4,30,0,2,30,2,2,30,3,5,189,1,2,
/* out0159_em-eta19-phi7*/	2,30,0,1,30,3,4,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	8,131,0,7,131,1,16,131,2,5,138,0,1,138,2,4,139,0,9,139,1,6,139,2,3,
/* out0164_em-eta4-phi8*/	6,120,1,10,120,2,6,121,0,2,121,1,1,131,0,8,131,2,4,
/* out0165_em-eta5-phi8*/	6,107,1,2,107,2,1,108,0,2,108,1,6,120,0,5,120,2,10,
/* out0166_em-eta6-phi8*/	3,95,1,4,107,2,9,108,0,8,
/* out0167_em-eta7-phi8*/	3,95,0,7,95,1,9,95,2,2,
/* out0168_em-eta8-phi8*/	4,82,1,6,82,2,1,95,0,7,226,1,8,
/* out0169_em-eta9-phi8*/	7,82,0,2,82,1,2,82,2,8,218,1,2,226,0,6,226,1,2,226,2,13,
/* out0170_em-eta10-phi8*/	9,67,5,4,68,5,2,69,1,4,70,1,7,82,0,2,82,2,3,218,1,12,218,2,2,219,0,2,
/* out0171_em-eta11-phi8*/	6,68,2,8,68,5,13,69,0,6,69,1,7,209,0,5,218,2,7,
/* out0172_em-eta12-phi8*/	8,50,4,10,51,1,5,68,2,8,68,3,3,69,0,1,208,1,3,209,0,7,209,2,1,
/* out0173_em-eta13-phi8*/	8,50,1,5,50,2,5,51,0,6,51,1,7,199,0,3,199,1,3,208,2,1,209,2,1,
/* out0174_em-eta14-phi8*/	7,50,0,8,50,1,3,50,2,5,50,3,4,199,0,5,199,1,1,199,2,2,
/* out0175_em-eta15-phi8*/	5,30,4,6,30,5,5,50,0,3,50,3,2,199,2,6,
/* out0176_em-eta16-phi8*/	5,30,5,4,31,0,8,31,4,2,189,0,2,189,2,5,
/* out0177_em-eta17-phi8*/	5,30,2,2,31,0,1,31,4,8,189,0,5,189,1,2,
/* out0178_em-eta18-phi8*/	5,30,2,2,30,3,2,31,3,3,31,4,2,189,1,1,
/* out0179_em-eta19-phi8*/	2,30,3,5,31,3,3,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	4,132,1,2,139,0,2,139,1,1,139,2,4,
/* out0183_em-eta3-phi9*/	7,131,2,5,132,0,15,132,1,12,132,2,2,139,0,5,139,1,9,139,2,9,
/* out0184_em-eta4-phi9*/	5,121,0,7,121,1,15,121,2,7,131,2,2,132,0,1,
/* out0185_em-eta5-phi9*/	6,108,1,10,108,2,5,109,0,1,109,1,1,121,0,7,121,2,2,
/* out0186_em-eta6-phi9*/	4,95,1,1,96,1,3,108,0,6,108,2,10,
/* out0187_em-eta7-phi9*/	4,83,1,1,95,1,2,95,2,10,96,0,5,
/* out0188_em-eta8-phi9*/	6,82,2,1,83,0,3,83,1,7,95,2,4,226,1,3,227,0,10,
/* out0189_em-eta9-phi9*/	9,69,4,5,82,2,3,83,0,8,219,0,6,219,1,5,226,1,2,226,2,3,227,0,2,227,2,3,
/* out0190_em-eta10-phi9*/	9,69,1,1,69,2,1,69,4,11,69,5,4,70,0,14,70,1,9,219,0,8,219,1,1,219,2,6,
/* out0191_em-eta11-phi9*/	8,69,0,5,69,1,4,69,2,15,69,3,6,70,4,2,209,0,2,209,1,9,219,2,2,
/* out0192_em-eta12-phi9*/	7,50,4,6,50,5,13,69,0,4,69,3,6,209,0,2,209,1,2,209,2,7,
/* out0193_em-eta13-phi9*/	7,50,2,1,50,5,1,51,0,10,51,4,10,51,5,2,199,1,5,209,2,4,
/* out0194_em-eta14-phi9*/	6,50,2,5,50,3,4,51,3,6,51,4,5,199,1,6,199,2,2,
/* out0195_em-eta15-phi9*/	7,30,5,5,31,5,1,32,1,1,50,3,6,51,3,3,190,0,1,199,2,5,
/* out0196_em-eta16-phi9*/	5,30,5,2,31,4,1,31,5,11,189,0,3,190,0,3,
/* out0197_em-eta17-phi9*/	6,31,2,4,31,3,1,31,4,3,31,5,3,189,0,6,190,0,2,
/* out0198_em-eta18-phi9*/	3,31,2,3,31,3,6,189,1,1,
/* out0199_em-eta19-phi9*/	2,13,4,3,31,3,3,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	1,132,1,1,
/* out0203_em-eta3-phi10*/	6,122,1,9,132,1,1,132,2,14,133,0,15,133,1,15,133,2,14,
/* out0204_em-eta4-phi10*/	5,109,1,3,121,2,6,122,0,15,122,1,5,122,2,1,
/* out0205_em-eta5-phi10*/	4,109,0,10,109,1,11,109,2,4,121,2,1,
/* out0206_em-eta6-phi10*/	5,96,1,12,96,2,3,108,2,1,109,0,5,109,2,1,
/* out0207_em-eta7-phi10*/	4,83,1,1,96,0,11,96,1,1,96,2,6,
/* out0208_em-eta8-phi10*/	5,83,1,7,83,2,7,220,0,1,227,0,4,227,2,6,
/* out0209_em-eta9-phi10*/	7,69,5,1,71,1,1,83,0,5,83,2,6,219,1,6,220,0,7,227,2,7,
/* out0210_em-eta10-phi10*/	10,69,5,11,70,0,2,70,2,3,70,4,5,70,5,15,71,0,1,210,0,3,219,1,4,219,2,7,220,0,1,
/* out0211_em-eta11-phi10*/	10,52,4,1,53,1,1,69,3,1,70,2,9,70,3,12,70,4,9,70,5,1,209,1,3,210,0,8,219,2,1,
/* out0212_em-eta12-phi10*/	12,50,5,2,51,5,4,52,1,7,53,1,7,69,3,3,70,3,4,200,0,2,200,1,1,209,1,2,209,2,3,210,0,1,210,2,1,
/* out0213_em-eta13-phi10*/	6,51,2,8,51,4,1,51,5,10,52,0,2,52,1,2,200,0,9,
/* out0214_em-eta14-phi10*/	7,32,4,4,33,1,1,51,2,8,51,3,6,199,1,1,200,0,4,200,2,2,
/* out0215_em-eta15-phi10*/	5,32,1,4,33,1,11,51,3,1,190,0,4,190,1,3,
/* out0216_em-eta16-phi10*/	5,31,2,1,31,5,1,32,0,2,32,1,9,190,0,5,
/* out0217_em-eta17-phi10*/	5,14,5,1,31,2,6,32,0,5,190,0,1,190,2,3,
/* out0218_em-eta18-phi10*/	4,13,4,2,13,5,11,31,2,2,190,2,1,
/* out0219_em-eta19-phi10*/	1,13,4,6,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	6,122,1,2,122,2,3,123,2,2,133,0,1,133,1,1,133,2,2,
/* out0224_em-eta4-phi11*/	6,109,1,1,110,0,2,110,1,12,122,0,1,122,2,12,123,2,3,
/* out0225_em-eta5-phi11*/	3,97,1,5,109,2,10,110,0,10,
/* out0226_em-eta6-phi11*/	4,96,2,3,97,0,10,97,1,7,109,2,1,
/* out0227_em-eta7-phi11*/	3,84,1,11,96,2,4,97,0,2,
/* out0228_em-eta8-phi11*/	5,83,2,2,84,0,12,84,1,1,220,0,1,220,1,5,
/* out0229_em-eta9-phi11*/	5,71,1,10,83,2,1,220,0,6,220,1,7,220,2,5,
/* out0230_em-eta10-phi11*/	6,70,2,1,71,0,9,71,1,1,210,0,1,210,1,8,220,2,7,
/* out0231_em-eta11-phi11*/	9,52,4,15,52,5,4,53,0,1,53,1,2,70,2,3,71,0,2,210,0,3,210,1,4,210,2,6,
/* out0232_em-eta12-phi11*/	6,52,1,3,52,2,8,53,0,11,53,1,6,200,1,5,210,2,5,
/* out0233_em-eta13-phi11*/	7,52,0,12,52,1,4,52,2,4,52,3,4,200,0,1,200,1,6,200,2,2,
/* out0234_em-eta14-phi11*/	6,32,4,12,32,5,4,33,0,1,33,1,1,52,0,2,200,2,8,
/* out0235_em-eta15-phi11*/	4,32,2,3,33,0,11,33,1,3,190,1,6,
/* out0236_em-eta16-phi11*/	6,32,0,1,32,1,2,32,2,9,32,3,1,190,1,3,190,2,3,
/* out0237_em-eta17-phi11*/	4,14,5,2,32,0,8,32,3,3,190,2,4,
/* out0238_em-eta18-phi11*/	5,13,5,4,14,0,6,14,4,4,14,5,9,190,2,1,
/* out0239_em-eta19-phi11*/	4,13,4,5,13,5,1,14,0,6,14,1,2,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	5,111,1,5,123,1,15,123,2,7,124,0,12,124,2,2,
/* out0244_em-eta4-phi12*/	7,98,1,1,110,1,4,110,2,10,111,0,8,111,1,4,123,1,1,123,2,4,
/* out0245_em-eta5-phi12*/	6,97,1,3,97,2,2,98,0,4,98,1,6,110,0,4,110,2,6,
/* out0246_em-eta6-phi12*/	5,85,1,3,97,0,3,97,1,1,97,2,14,98,0,1,
/* out0247_em-eta7-phi12*/	5,84,1,4,84,2,7,85,0,3,85,1,1,97,0,1,
/* out0248_em-eta8-phi12*/	4,72,1,2,84,0,4,84,2,9,221,0,8,
/* out0249_em-eta9-phi12*/	9,71,1,4,71,2,7,72,0,1,211,0,3,211,1,3,220,1,4,220,2,3,221,0,5,221,2,4,
/* out0250_em-eta10-phi12*/	7,55,1,1,71,0,2,71,2,7,210,1,1,211,0,12,211,2,1,220,2,1,
/* out0251_em-eta11-phi12*/	12,52,5,12,53,0,1,53,5,10,54,1,2,55,1,2,71,0,2,201,0,3,201,1,2,210,1,3,210,2,3,211,0,1,211,2,1,
/* out0252_em-eta12-phi12*/	9,52,2,1,53,0,3,53,2,2,53,3,3,53,4,15,53,5,5,200,1,1,201,0,9,210,2,1,
/* out0253_em-eta13-phi12*/	9,52,2,3,52,3,10,53,3,9,53,4,1,191,0,1,200,1,3,200,2,2,201,0,2,201,2,1,
/* out0254_em-eta14-phi12*/	6,32,5,12,33,0,1,33,5,5,52,3,2,191,0,5,200,2,2,
/* out0255_em-eta15-phi12*/	5,33,0,3,33,4,10,33,5,2,190,1,2,191,0,4,
/* out0256_em-eta16-phi12*/	8,32,2,4,32,3,1,33,3,3,33,4,6,181,1,1,190,1,2,190,2,2,191,0,1,
/* out0257_em-eta17-phi12*/	5,14,2,1,32,3,10,33,3,1,181,1,3,190,2,2,
/* out0258_em-eta18-phi12*/	5,14,2,7,14,3,1,14,4,6,14,5,4,181,1,1,
/* out0259_em-eta19-phi12*/	5,13,1,4,13,3,4,14,0,4,14,1,8,14,4,5,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	1,112,1,1,
/* out0263_em-eta3-phi13*/	6,111,1,5,111,2,4,112,0,6,112,1,8,124,0,4,124,2,14,
/* out0264_em-eta4-phi13*/	8,98,1,3,98,2,1,99,0,2,99,1,4,111,0,8,111,1,2,111,2,12,112,0,1,
/* out0265_em-eta5-phi13*/	4,98,0,6,98,1,6,98,2,13,99,0,1,
/* out0266_em-eta6-phi13*/	5,85,1,11,85,2,4,86,1,1,98,0,5,98,2,1,
/* out0267_em-eta7-phi13*/	4,72,1,1,85,0,13,85,1,1,85,2,3,
/* out0268_em-eta8-phi13*/	6,72,0,1,72,1,13,72,2,1,212,0,2,221,0,3,221,2,5,
/* out0269_em-eta9-phi13*/	6,54,4,1,71,2,1,72,0,11,211,1,7,212,0,6,221,2,7,
/* out0270_em-eta10-phi13*/	7,54,4,15,54,5,3,55,0,7,55,1,10,71,2,1,211,1,6,211,2,9,
/* out0271_em-eta11-phi13*/	9,53,5,1,54,0,5,54,1,14,54,2,7,55,0,2,55,1,3,201,1,8,202,0,1,211,2,4,
/* out0272_em-eta12-phi13*/	6,34,4,7,53,2,13,54,0,7,201,0,2,201,1,3,201,2,5,
/* out0273_em-eta13-phi13*/	7,34,4,3,35,0,1,35,1,15,53,2,1,53,3,4,191,1,4,201,2,5,
/* out0274_em-eta14-phi13*/	5,33,5,5,34,0,2,34,1,13,191,0,2,191,1,5,
/* out0275_em-eta15-phi13*/	5,33,2,11,33,5,4,34,0,1,191,0,3,191,2,4,
/* out0276_em-eta16-phi13*/	7,15,4,1,16,1,1,33,2,4,33,3,8,181,1,1,181,2,3,191,2,2,
/* out0277_em-eta17-phi13*/	7,14,2,1,15,1,1,16,1,5,32,3,1,33,3,4,181,1,5,181,2,1,
/* out0278_em-eta18-phi13*/	4,14,2,7,14,3,5,15,1,2,181,1,1,
/* out0279_em-eta19-phi13*/	5,13,1,10,13,3,10,14,1,5,14,3,6,14,4,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	5,112,1,2,112,2,1,113,0,4,113,1,1,113,2,2,
/* out0283_em-eta3-phi14*/	8,100,0,1,100,1,5,112,0,8,112,1,5,112,2,15,113,0,9,113,1,9,113,2,5,
/* out0284_em-eta4-phi14*/	5,99,0,5,99,1,12,99,2,12,100,0,1,112,0,1,
/* out0285_em-eta5-phi14*/	5,86,1,13,86,2,2,98,2,1,99,0,8,99,2,1,
/* out0286_em-eta6-phi14*/	5,73,1,1,85,2,4,86,0,13,86,1,2,86,2,1,
/* out0287_em-eta7-phi14*/	3,73,0,3,73,1,9,85,2,5,
/* out0288_em-eta8-phi14*/	7,56,1,1,72,2,10,73,0,4,212,0,1,212,1,10,213,0,1,213,1,1,
/* out0289_em-eta9-phi14*/	9,54,5,4,55,5,1,56,0,1,56,1,2,72,0,3,72,2,5,212,0,7,212,1,3,212,2,9,
/* out0290_em-eta10-phi14*/	9,54,5,9,55,0,6,55,2,1,55,4,8,55,5,15,202,0,6,202,1,7,211,2,1,212,2,2,
/* out0291_em-eta11-phi14*/	8,54,2,9,54,3,9,55,0,1,55,3,7,55,4,8,201,1,1,202,0,9,202,2,2,
/* out0292_em-eta12-phi14*/	9,34,4,5,34,5,13,54,0,4,54,3,6,192,0,4,192,1,1,201,1,2,201,2,4,202,2,1,
/* out0293_em-eta13-phi14*/	9,34,2,3,34,4,1,34,5,1,35,0,15,35,1,1,35,4,3,191,1,2,192,0,6,201,2,1,
/* out0294_em-eta14-phi14*/	6,34,0,4,34,1,3,34,2,10,34,3,3,191,1,5,191,2,2,
/* out0295_em-eta15-phi14*/	4,15,4,6,33,2,1,34,0,9,191,2,6,
/* out0296_em-eta16-phi14*/	5,15,4,8,16,0,1,16,1,5,181,2,5,191,2,1,
/* out0297_em-eta17-phi14*/	6,15,1,3,15,2,1,16,0,2,16,1,5,181,1,3,181,2,3,
/* out0298_em-eta18-phi14*/	2,15,0,1,15,1,8,
/* out0299_em-eta19-phi14*/	5,13,1,2,13,3,2,14,1,1,14,3,4,15,0,3,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	7,100,0,3,100,1,11,100,2,13,101,0,6,113,0,3,113,1,6,113,2,9,
/* out0304_em-eta4-phi15*/	5,87,1,14,87,2,2,99,2,3,100,0,11,100,2,2,
/* out0305_em-eta5-phi15*/	4,74,1,2,86,2,7,87,0,13,87,1,2,
/* out0306_em-eta6-phi15*/	6,73,1,2,73,2,2,74,0,3,74,1,6,86,0,3,86,2,6,
/* out0307_em-eta7-phi15*/	3,73,0,2,73,1,4,73,2,11,
/* out0308_em-eta8-phi15*/	8,56,1,7,73,0,7,73,2,1,203,1,1,212,1,2,213,0,14,213,1,14,213,2,14,
/* out0309_em-eta9-phi15*/	7,56,0,5,56,1,6,56,2,1,203,0,9,203,1,3,212,1,1,212,2,5,
/* out0310_em-eta10-phi15*/	6,36,4,6,55,2,11,56,0,6,202,1,9,202,2,2,203,0,4,
/* out0311_em-eta11-phi15*/	7,36,4,6,37,1,14,55,2,4,55,3,9,192,1,1,193,0,1,202,2,11,
/* out0312_em-eta12-phi15*/	9,34,5,2,35,2,1,35,5,12,36,0,1,36,1,10,37,1,1,54,3,1,192,0,1,192,1,10,
/* out0313_em-eta13-phi15*/	6,35,2,5,35,3,3,35,4,11,35,5,4,192,0,4,192,2,4,
/* out0314_em-eta14-phi15*/	9,34,2,3,34,3,8,35,3,7,35,4,2,182,0,1,182,1,3,191,2,1,192,0,1,192,2,2,
/* out0315_em-eta15-phi15*/	4,15,4,1,15,5,10,34,3,5,182,0,6,
/* out0316_em-eta16-phi15*/	4,15,5,4,16,0,9,181,2,1,182,0,4,
/* out0317_em-eta17-phi15*/	5,15,2,7,16,0,4,16,4,1,181,1,1,181,2,3,
/* out0318_em-eta18-phi15*/	4,15,0,3,15,1,2,15,2,4,15,3,1,
/* out0319_em-eta19-phi15*/	1,15,0,7,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	3,89,0,3,101,0,4,101,2,3,
/* out0323_em-eta3-phi16*/	7,88,1,13,88,2,6,89,0,3,89,2,1,100,2,1,101,0,6,101,2,13,
/* out0324_em-eta4-phi16*/	5,75,1,4,87,2,9,88,0,14,88,1,3,88,2,1,
/* out0325_em-eta5-phi16*/	6,74,1,4,74,2,4,75,0,4,75,1,5,87,0,3,87,2,5,
/* out0326_em-eta6-phi16*/	3,74,0,10,74,1,4,74,2,8,
/* out0327_em-eta7-phi16*/	3,57,1,12,73,2,2,74,0,3,
/* out0328_em-eta8-phi16*/	10,56,2,5,57,0,8,57,1,2,203,1,3,204,0,6,204,1,4,204,2,3,213,0,1,213,1,1,213,2,2,
/* out0329_em-eta9-phi16*/	8,38,1,1,56,0,1,56,2,10,203,0,2,203,1,9,203,2,7,204,0,2,204,1,1,
/* out0330_em-eta10-phi16*/	8,36,4,3,36,5,15,37,5,5,56,0,3,193,0,1,193,1,6,203,0,1,203,2,7,
/* out0331_em-eta11-phi16*/	8,36,2,8,36,4,1,36,5,1,37,0,16,37,1,1,37,4,7,193,0,11,193,1,2,
/* out0332_em-eta12-phi16*/	10,35,2,1,36,0,12,36,1,6,36,2,7,36,3,3,183,0,1,192,1,4,192,2,2,193,0,3,193,2,1,
/* out0333_em-eta13-phi16*/	6,17,4,11,18,1,1,35,2,9,36,0,2,183,0,2,192,2,7,
/* out0334_em-eta14-phi16*/	5,17,1,2,18,1,12,35,3,6,182,1,6,192,2,1,
/* out0335_em-eta15-phi16*/	6,15,5,2,16,5,9,17,1,5,182,0,2,182,1,3,182,2,2,
/* out0336_em-eta16-phi16*/	4,16,4,7,16,5,7,182,0,2,182,2,3,
/* out0337_em-eta17-phi16*/	5,15,2,2,16,3,1,16,4,8,182,0,1,182,2,1,
/* out0338_em-eta18-phi16*/	3,15,2,2,15,3,7,16,3,1,
/* out0339_em-eta19-phi16*/	2,15,0,2,15,3,3,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	1,89,0,2,
/* out0343_em-eta3-phi17*/	4,76,1,11,88,2,5,89,0,8,89,2,15,
/* out0344_em-eta4-phi17*/	6,75,1,5,75,2,8,76,0,8,76,1,5,88,0,2,88,2,4,
/* out0345_em-eta5-phi17*/	5,58,1,4,74,2,1,75,0,12,75,1,2,75,2,8,
/* out0346_em-eta6-phi17*/	3,58,0,5,58,1,12,74,2,3,
/* out0347_em-eta7-phi17*/	3,57,1,2,57,2,13,58,0,3,
/* out0348_em-eta8-phi17*/	7,38,1,4,57,0,8,57,2,3,194,1,1,204,0,6,204,1,4,204,2,9,
/* out0349_em-eta9-phi17*/	8,38,0,1,38,1,11,194,0,7,194,1,7,203,2,2,204,0,2,204,1,7,204,2,4,
/* out0350_em-eta10-phi17*/	5,37,2,5,37,5,8,38,0,7,193,1,6,194,0,9,
/* out0351_em-eta11-phi17*/	6,37,2,11,37,3,11,37,4,9,37,5,3,193,1,2,193,2,11,
/* out0352_em-eta12-phi17*/	8,17,4,1,17,5,6,36,0,1,36,2,1,36,3,13,37,3,5,183,1,7,193,2,4,
/* out0353_em-eta13-phi17*/	6,17,4,4,17,5,10,18,0,9,18,1,1,183,0,8,183,1,1,
/* out0354_em-eta14-phi17*/	6,17,1,2,17,2,7,18,0,7,18,1,2,182,1,3,183,0,5,
/* out0355_em-eta15-phi17*/	6,16,2,1,17,0,7,17,1,7,17,2,1,182,1,1,182,2,5,
/* out0356_em-eta16-phi17*/	3,16,2,13,17,0,1,182,2,5,
/* out0357_em-eta17-phi17*/	2,16,2,2,16,3,9,
/* out0358_em-eta18-phi17*/	2,15,3,4,16,3,5,
/* out0359_em-eta19-phi17*/	1,15,3,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	1,77,0,2,
/* out0363_em-eta3-phi18*/	4,60,1,5,76,2,11,77,0,14,77,2,9,
/* out0364_em-eta4-phi18*/	6,59,1,8,59,2,5,60,0,2,60,1,4,76,0,8,76,2,5,
/* out0365_em-eta5-phi18*/	5,40,1,1,58,2,4,59,0,12,59,1,8,59,2,2,
/* out0366_em-eta6-phi18*/	3,40,1,3,58,0,5,58,2,12,
/* out0367_em-eta7-phi18*/	3,39,1,13,39,2,2,58,0,3,
/* out0368_em-eta8-phi18*/	7,38,2,4,39,0,8,39,1,3,194,1,1,195,0,9,195,1,4,195,2,6,
/* out0369_em-eta9-phi18*/	8,38,0,1,38,2,11,185,0,2,194,1,7,194,2,7,195,0,4,195,1,7,195,2,2,
/* out0370_em-eta10-phi18*/	5,19,4,5,19,5,8,38,0,7,184,1,6,194,2,9,
/* out0371_em-eta11-phi18*/	6,19,4,11,19,5,3,20,0,9,20,1,11,184,0,11,184,1,2,
/* out0372_em-eta12-phi18*/	8,18,2,1,18,5,6,19,0,1,19,1,13,19,2,1,20,1,5,183,1,7,184,0,4,
/* out0373_em-eta13-phi18*/	6,18,2,4,18,3,1,18,4,9,18,5,10,183,1,1,183,2,8,
/* out0374_em-eta14-phi18*/	6,17,2,7,17,3,2,18,3,2,18,4,7,177,1,3,183,2,5,
/* out0375_em-eta15-phi18*/	6,0,4,1,17,0,7,17,2,1,17,3,7,177,0,5,177,1,1,
/* out0376_em-eta16-phi18*/	3,0,4,13,17,0,1,177,0,5,
/* out0377_em-eta17-phi18*/	2,0,4,2,1,1,9,
/* out0378_em-eta18-phi18*/	2,0,1,4,1,1,5,
/* out0379_em-eta19-phi18*/	1,0,1,1,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	2,61,0,7,77,2,2,
/* out0383_em-eta3-phi19*/	6,42,1,1,60,1,6,60,2,13,61,0,8,61,2,12,77,2,5,
/* out0384_em-eta4-phi19*/	5,41,1,9,59,2,4,60,0,14,60,1,1,60,2,3,
/* out0385_em-eta5-phi19*/	6,40,1,4,40,2,4,41,0,3,41,1,5,59,0,4,59,2,5,
/* out0386_em-eta6-phi19*/	3,40,0,10,40,1,8,40,2,4,
/* out0387_em-eta7-phi19*/	3,22,1,2,39,2,12,40,0,3,
/* out0388_em-eta8-phi19*/	10,21,1,5,39,0,8,39,2,2,185,1,3,186,0,2,186,1,1,186,2,1,195,0,3,195,1,4,195,2,6,
/* out0389_em-eta9-phi19*/	8,21,0,1,21,1,10,38,2,1,185,0,7,185,1,9,185,2,2,195,1,1,195,2,2,
/* out0390_em-eta10-phi19*/	8,19,5,5,20,2,3,20,5,15,21,0,3,184,1,6,184,2,1,185,0,7,185,2,1,
/* out0391_em-eta11-phi19*/	8,19,2,8,20,0,7,20,2,1,20,3,1,20,4,16,20,5,1,184,1,2,184,2,11,
/* out0392_em-eta12-phi19*/	10,2,4,1,19,0,12,19,1,3,19,2,7,19,3,6,178,0,2,178,1,4,183,2,1,184,0,1,184,2,3,
/* out0393_em-eta13-phi19*/	6,2,4,9,18,2,11,18,3,1,19,0,2,178,0,7,183,2,2,
/* out0394_em-eta14-phi19*/	5,3,1,6,17,3,2,18,3,12,177,1,6,178,0,1,
/* out0395_em-eta15-phi19*/	6,0,5,9,1,5,2,17,3,5,177,0,2,177,1,3,177,2,2,
/* out0396_em-eta16-phi19*/	4,0,5,7,1,0,7,177,0,3,177,2,2,
/* out0397_em-eta17-phi19*/	5,0,2,2,1,0,8,1,1,1,177,0,1,177,2,1,
/* out0398_em-eta18-phi19*/	3,0,1,7,0,2,2,1,1,1,
/* out0399_em-eta19-phi19*/	2,0,0,2,0,1,3,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	8,42,0,3,42,1,13,42,2,11,43,0,9,43,1,6,43,2,3,61,0,1,61,2,4,
/* out0404_em-eta4-phi20*/	5,24,1,3,41,1,2,41,2,14,42,0,11,42,1,2,
/* out0405_em-eta5-phi20*/	4,23,1,7,40,2,2,41,0,13,41,2,2,
/* out0406_em-eta6-phi20*/	6,22,1,2,22,2,2,23,0,3,23,1,6,40,0,3,40,2,6,
/* out0407_em-eta7-phi20*/	3,22,0,2,22,1,11,22,2,4,
/* out0408_em-eta8-phi20*/	8,21,2,7,22,0,7,22,1,1,180,1,2,185,1,1,186,0,14,186,1,14,186,2,14,
/* out0409_em-eta9-phi20*/	7,21,0,5,21,1,1,21,2,6,180,0,5,180,1,1,185,1,3,185,2,9,
/* out0410_em-eta10-phi20*/	6,4,4,11,20,2,6,21,0,6,179,0,2,179,1,9,185,2,4,
/* out0411_em-eta11-phi20*/	7,4,4,4,5,1,9,20,2,6,20,3,14,178,1,1,179,0,11,184,2,1,
/* out0412_em-eta12-phi20*/	9,2,4,1,2,5,12,3,5,2,4,1,1,19,0,1,19,3,10,20,3,1,178,1,10,178,2,1,
/* out0413_em-eta13-phi20*/	6,2,4,5,2,5,4,3,0,11,3,1,3,178,0,4,178,2,4,
/* out0414_em-eta14-phi20*/	9,2,1,8,2,2,3,3,0,2,3,1,7,173,0,1,177,1,3,177,2,1,178,0,2,178,2,1,
/* out0415_em-eta15-phi20*/	4,1,2,1,1,5,10,2,1,5,177,2,6,
/* out0416_em-eta16-phi20*/	4,1,4,9,1,5,4,172,1,1,177,2,4,
/* out0417_em-eta17-phi20*/	4,0,2,7,1,0,1,1,4,4,172,1,4,
/* out0418_em-eta18-phi20*/	4,0,0,3,0,1,1,0,2,4,0,3,2,
/* out0419_em-eta19-phi20*/	1,0,0,7,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	5,25,1,1,25,2,2,43,0,2,43,1,1,43,2,4,
/* out0423_em-eta3-phi21*/	8,25,0,8,25,1,15,25,2,5,42,0,1,42,2,5,43,0,5,43,1,9,43,2,9,
/* out0424_em-eta4-phi21*/	5,24,0,5,24,1,12,24,2,12,25,0,1,42,0,1,
/* out0425_em-eta5-phi21*/	5,8,1,1,23,1,2,23,2,13,24,0,8,24,1,1,
/* out0426_em-eta6-phi21*/	5,7,1,4,22,2,1,23,0,13,23,1,1,23,2,2,
/* out0427_em-eta7-phi21*/	3,7,1,5,22,0,3,22,2,9,
/* out0428_em-eta8-phi21*/	7,6,1,10,21,2,1,22,0,4,180,1,10,180,2,1,186,1,1,186,2,1,
/* out0429_em-eta9-phi21*/	9,4,5,1,5,5,4,6,0,3,6,1,5,21,0,1,21,2,2,180,0,9,180,1,3,180,2,7,
/* out0430_em-eta10-phi21*/	9,4,4,1,4,5,15,5,0,8,5,4,6,5,5,9,175,0,1,179,1,7,179,2,6,180,0,2,
/* out0431_em-eta11-phi21*/	8,4,1,9,4,2,9,5,0,8,5,1,7,5,4,1,174,1,1,179,0,2,179,2,9,
/* out0432_em-eta12-phi21*/	9,3,2,5,3,5,13,4,0,4,4,1,6,174,0,4,174,1,2,178,1,1,178,2,4,179,0,1,
/* out0433_em-eta13-phi21*/	9,2,2,3,3,0,3,3,2,1,3,3,1,3,4,15,3,5,1,173,1,2,174,0,1,178,2,6,
/* out0434_em-eta14-phi21*/	6,2,0,4,2,1,3,2,2,10,2,3,3,173,0,2,173,1,5,
/* out0435_em-eta15-phi21*/	3,1,2,6,2,0,9,173,0,6,
/* out0436_em-eta16-phi21*/	6,1,2,8,1,3,5,1,4,1,172,1,2,172,2,3,173,0,1,
/* out0437_em-eta17-phi21*/	6,0,2,1,0,3,3,1,3,5,1,4,2,172,1,5,172,2,1,
/* out0438_em-eta18-phi21*/	2,0,0,1,0,3,8,
/* out0439_em-eta19-phi21*/	1,0,0,3,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	1,25,2,1,
/* out0443_em-eta3-phi22*/	7,9,1,4,9,2,5,10,0,15,10,1,15,10,2,14,25,0,6,25,2,8,
/* out0444_em-eta4-phi22*/	8,8,1,1,8,2,3,9,0,8,9,1,12,9,2,2,24,0,2,24,2,4,25,0,1,
/* out0445_em-eta5-phi22*/	4,8,0,6,8,1,13,8,2,6,24,0,1,
/* out0446_em-eta6-phi22*/	5,7,1,4,7,2,11,8,0,5,8,1,1,23,2,1,
/* out0447_em-eta7-phi22*/	4,6,2,1,7,0,13,7,1,3,7,2,1,
/* out0448_em-eta8-phi22*/	5,6,0,1,6,1,1,6,2,13,176,0,8,180,2,2,
/* out0449_em-eta9-phi22*/	6,5,2,1,6,0,11,175,1,7,176,0,4,176,2,3,180,2,6,
/* out0450_em-eta10-phi22*/	6,5,2,15,5,3,10,5,4,7,5,5,3,175,0,9,175,1,6,
/* out0451_em-eta11-phi22*/	8,4,0,5,4,2,7,4,3,14,5,3,3,5,4,2,174,1,8,175,0,4,179,2,1,
/* out0452_em-eta12-phi22*/	5,3,2,7,4,0,7,174,0,5,174,1,3,174,2,2,
/* out0453_em-eta13-phi22*/	5,3,2,3,3,3,15,3,4,1,173,1,4,174,0,5,
/* out0454_em-eta14-phi22*/	4,2,0,2,2,3,13,173,1,5,173,2,2,
/* out0455_em-eta15-phi22*/	3,2,0,1,173,0,4,173,2,3,
/* out0456_em-eta16-phi22*/	4,1,2,1,1,3,1,172,2,4,173,0,2,
/* out0457_em-eta17-phi22*/	4,0,3,1,1,3,5,172,1,2,172,2,4,
/* out0458_em-eta18-phi22*/	2,0,3,2,172,1,1,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	4,9,2,5,10,0,1,10,1,1,10,2,2,
/* out0464_em-eta4-phi23*/	3,8,2,1,9,0,8,9,2,4,
/* out0465_em-eta5-phi23*/	2,8,0,4,8,2,6,
/* out0466_em-eta6-phi23*/	2,7,2,3,8,0,1,
/* out0467_em-eta7-phi23*/	2,7,0,3,7,2,1,
/* out0468_em-eta8-phi23*/	3,6,2,2,176,0,4,176,2,4,
/* out0469_em-eta9-phi23*/	4,6,0,1,175,1,3,175,2,3,176,2,9,
/* out0470_em-eta10-phi23*/	3,5,3,1,175,0,1,175,2,12,
/* out0471_em-eta11-phi23*/	6,4,3,2,5,3,2,174,1,2,174,2,3,175,0,1,175,2,1,
/* out0472_em-eta12-phi23*/	1,174,2,9,
/* out0473_em-eta13-phi23*/	3,173,2,1,174,0,1,174,2,2,
/* out0474_em-eta14-phi23*/	1,173,2,5,
/* out0475_em-eta15-phi23*/	1,173,2,4,
/* out0476_em-eta16-phi23*/	2,172,2,1,173,2,1,
/* out0477_em-eta17-phi23*/	1,172,2,3,
/* out0478_em-eta18-phi23*/	1,172,1,1,
/* out0479_em-eta19-phi23*/	0
};