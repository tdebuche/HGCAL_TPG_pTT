parameter integer matrixH [0:2516] = {
/* num inputs = 174(in0-in173) */
/* num outputs = 560(out0-out559) */
//* max inputs per outputs = 5 */
//* total number of input in adders 978 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	1, 0, 1, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	0, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	1, 3, 1, 
/* out0033_had-eta13-phi1*/	0, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	1, 1, 1, 
/* out0036_had-eta16-phi1*/	1, 1, 1, 
/* out0037_had-eta17-phi1*/	0, 
/* out0038_had-eta18-phi1*/	1, 0, 2, 
/* out0039_had-eta19-phi1*/	1, 0, 1, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	1, 27, 4, 
/* out0045_had-eta5-phi2*/	2, 26, 1, 27, 4, 
/* out0046_had-eta6-phi2*/	1, 26, 6, 
/* out0047_had-eta7-phi2*/	2, 25, 3, 26, 1, 
/* out0048_had-eta8-phi2*/	1, 25, 5, 
/* out0049_had-eta9-phi2*/	1, 24, 3, 
/* out0050_had-eta10-phi2*/	1, 24, 3, 
/* out0051_had-eta11-phi2*/	2, 3, 2, 24, 1, 
/* out0052_had-eta12-phi2*/	1, 3, 2, 
/* out0053_had-eta13-phi2*/	1, 3, 2, 
/* out0054_had-eta14-phi2*/	1, 1, 2, 
/* out0055_had-eta15-phi2*/	1, 1, 1, 
/* out0056_had-eta16-phi2*/	1, 1, 1, 
/* out0057_had-eta17-phi2*/	1, 1, 1, 
/* out0058_had-eta18-phi2*/	1, 0, 2, 
/* out0059_had-eta19-phi2*/	1, 0, 2, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 118, 4, 
/* out0062_had-eta2-phi3*/	1, 118, 4, 
/* out0063_had-eta3-phi3*/	3, 35, 1, 36, 7, 117, 5, 
/* out0064_had-eta4-phi3*/	4, 27, 4, 35, 5, 116, 1, 117, 3, 
/* out0065_had-eta5-phi3*/	4, 26, 1, 27, 4, 34, 3, 116, 4, 
/* out0066_had-eta6-phi3*/	5, 26, 6, 33, 1, 34, 1, 115, 1, 116, 3, 
/* out0067_had-eta7-phi3*/	4, 25, 3, 26, 1, 33, 2, 115, 3, 
/* out0068_had-eta8-phi3*/	2, 25, 5, 115, 3, 
/* out0069_had-eta9-phi3*/	4, 24, 3, 32, 1, 114, 3, 115, 1, 
/* out0070_had-eta10-phi3*/	2, 24, 4, 114, 5, 
/* out0071_had-eta11-phi3*/	2, 3, 2, 24, 1, 
/* out0072_had-eta12-phi3*/	1, 3, 3, 
/* out0073_had-eta13-phi3*/	1, 3, 2, 
/* out0074_had-eta14-phi3*/	1, 1, 2, 
/* out0075_had-eta15-phi3*/	1, 1, 1, 
/* out0076_had-eta16-phi3*/	1, 1, 1, 
/* out0077_had-eta17-phi3*/	1, 1, 1, 
/* out0078_had-eta18-phi3*/	1, 0, 2, 
/* out0079_had-eta19-phi3*/	1, 0, 2, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 118, 4, 
/* out0082_had-eta2-phi4*/	1, 118, 4, 
/* out0083_had-eta3-phi4*/	4, 35, 2, 36, 9, 46, 5, 117, 5, 
/* out0084_had-eta4-phi4*/	5, 35, 8, 45, 2, 46, 1, 116, 1, 117, 3, 
/* out0085_had-eta5-phi4*/	2, 34, 8, 116, 4, 
/* out0086_had-eta6-phi4*/	4, 33, 4, 34, 3, 115, 1, 116, 3, 
/* out0087_had-eta7-phi4*/	2, 33, 6, 115, 3, 
/* out0088_had-eta8-phi4*/	2, 32, 5, 115, 3, 
/* out0089_had-eta9-phi4*/	3, 32, 4, 114, 3, 115, 1, 
/* out0090_had-eta10-phi4*/	3, 9, 3, 24, 1, 114, 5, 
/* out0091_had-eta11-phi4*/	1, 9, 3, 
/* out0092_had-eta12-phi4*/	3, 3, 1, 8, 1, 9, 1, 
/* out0093_had-eta13-phi4*/	2, 3, 1, 8, 2, 
/* out0094_had-eta14-phi4*/	2, 1, 1, 8, 1, 
/* out0095_had-eta15-phi4*/	1, 1, 1, 
/* out0096_had-eta16-phi4*/	1, 1, 1, 
/* out0097_had-eta17-phi4*/	2, 1, 1, 2, 1, 
/* out0098_had-eta18-phi4*/	1, 0, 2, 
/* out0099_had-eta19-phi4*/	1, 0, 1, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 123, 4, 
/* out0102_had-eta2-phi5*/	2, 56, 2, 123, 4, 
/* out0103_had-eta3-phi5*/	4, 46, 9, 55, 1, 56, 4, 122, 5, 
/* out0104_had-eta4-phi5*/	5, 45, 9, 46, 1, 55, 1, 121, 1, 122, 3, 
/* out0105_had-eta5-phi5*/	4, 34, 1, 44, 4, 45, 4, 121, 4, 
/* out0106_had-eta6-phi5*/	4, 33, 1, 44, 6, 120, 1, 121, 3, 
/* out0107_had-eta7-phi5*/	3, 33, 2, 43, 4, 120, 3, 
/* out0108_had-eta8-phi5*/	3, 32, 3, 43, 2, 120, 3, 
/* out0109_had-eta9-phi5*/	4, 32, 3, 42, 1, 119, 3, 120, 1, 
/* out0110_had-eta10-phi5*/	2, 9, 3, 119, 5, 
/* out0111_had-eta11-phi5*/	1, 9, 3, 
/* out0112_had-eta12-phi5*/	2, 8, 1, 9, 1, 
/* out0113_had-eta13-phi5*/	1, 8, 2, 
/* out0114_had-eta14-phi5*/	1, 8, 2, 
/* out0115_had-eta15-phi5*/	1, 8, 1, 
/* out0116_had-eta16-phi5*/	1, 2, 1, 
/* out0117_had-eta17-phi5*/	1, 2, 1, 
/* out0118_had-eta18-phi5*/	1, 2, 1, 
/* out0119_had-eta19-phi5*/	1, 0, 1, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 123, 4, 
/* out0122_had-eta2-phi6*/	3, 56, 5, 96, 2, 123, 4, 
/* out0123_had-eta3-phi6*/	4, 55, 8, 56, 5, 96, 3, 122, 5, 
/* out0124_had-eta4-phi6*/	5, 45, 1, 54, 5, 55, 6, 121, 1, 122, 3, 
/* out0125_had-eta5-phi6*/	4, 44, 2, 53, 1, 54, 6, 121, 4, 
/* out0126_had-eta6-phi6*/	5, 43, 1, 44, 4, 53, 3, 120, 1, 121, 3, 
/* out0127_had-eta7-phi6*/	2, 43, 6, 120, 3, 
/* out0128_had-eta8-phi6*/	3, 42, 2, 43, 3, 120, 3, 
/* out0129_had-eta9-phi6*/	3, 42, 4, 119, 3, 120, 1, 
/* out0130_had-eta10-phi6*/	3, 9, 1, 42, 2, 119, 5, 
/* out0131_had-eta11-phi6*/	2, 9, 1, 10, 2, 
/* out0132_had-eta12-phi6*/	2, 8, 1, 10, 1, 
/* out0133_had-eta13-phi6*/	1, 8, 2, 
/* out0134_had-eta14-phi6*/	1, 8, 2, 
/* out0135_had-eta15-phi6*/	1, 2, 1, 
/* out0136_had-eta16-phi6*/	1, 2, 1, 
/* out0137_had-eta17-phi6*/	1, 2, 1, 
/* out0138_had-eta18-phi6*/	1, 2, 1, 
/* out0139_had-eta19-phi6*/	1, 2, 1, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 128, 4, 
/* out0142_had-eta2-phi7*/	3, 96, 4, 97, 1, 128, 4, 
/* out0143_had-eta3-phi7*/	4, 95, 5, 96, 7, 97, 3, 127, 5, 
/* out0144_had-eta4-phi7*/	5, 54, 2, 94, 1, 95, 8, 126, 1, 127, 3, 
/* out0145_had-eta5-phi7*/	4, 53, 2, 54, 3, 94, 4, 126, 4, 
/* out0146_had-eta6-phi7*/	3, 53, 7, 125, 1, 126, 3, 
/* out0147_had-eta7-phi7*/	3, 52, 4, 53, 2, 125, 3, 
/* out0148_had-eta8-phi7*/	3, 42, 1, 52, 4, 125, 3, 
/* out0149_had-eta9-phi7*/	3, 42, 4, 124, 3, 125, 1, 
/* out0150_had-eta10-phi7*/	3, 10, 2, 42, 2, 124, 5, 
/* out0151_had-eta11-phi7*/	1, 10, 3, 
/* out0152_had-eta12-phi7*/	1, 10, 2, 
/* out0153_had-eta13-phi7*/	2, 8, 1, 14, 1, 
/* out0154_had-eta14-phi7*/	1, 14, 1, 
/* out0155_had-eta15-phi7*/	1, 2, 1, 
/* out0156_had-eta16-phi7*/	1, 2, 1, 
/* out0157_had-eta17-phi7*/	1, 2, 1, 
/* out0158_had-eta18-phi7*/	1, 2, 1, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 128, 4, 
/* out0162_had-eta2-phi8*/	1, 128, 4, 
/* out0163_had-eta3-phi8*/	4, 95, 1, 97, 12, 104, 3, 127, 5, 
/* out0164_had-eta4-phi8*/	5, 94, 3, 95, 2, 104, 5, 126, 1, 127, 3, 
/* out0165_had-eta5-phi8*/	2, 94, 8, 126, 4, 
/* out0166_had-eta6-phi8*/	4, 53, 1, 102, 6, 125, 1, 126, 3, 
/* out0167_had-eta7-phi8*/	3, 52, 4, 102, 1, 125, 3, 
/* out0168_had-eta8-phi8*/	3, 52, 4, 62, 1, 125, 3, 
/* out0169_had-eta9-phi8*/	3, 62, 4, 124, 3, 125, 1, 
/* out0170_had-eta10-phi8*/	3, 10, 1, 62, 3, 124, 5, 
/* out0171_had-eta11-phi8*/	1, 10, 3, 
/* out0172_had-eta12-phi8*/	1, 10, 2, 
/* out0173_had-eta13-phi8*/	1, 14, 2, 
/* out0174_had-eta14-phi8*/	1, 14, 2, 
/* out0175_had-eta15-phi8*/	1, 14, 1, 
/* out0176_had-eta16-phi8*/	1, 2, 1, 
/* out0177_had-eta17-phi8*/	1, 2, 1, 
/* out0178_had-eta18-phi8*/	1, 2, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 133, 4, 
/* out0182_had-eta2-phi9*/	1, 133, 4, 
/* out0183_had-eta3-phi9*/	4, 104, 3, 105, 1, 106, 12, 132, 5, 
/* out0184_had-eta4-phi9*/	5, 103, 3, 104, 5, 105, 2, 131, 1, 132, 3, 
/* out0185_had-eta5-phi9*/	3, 102, 1, 103, 8, 131, 4, 
/* out0186_had-eta6-phi9*/	4, 64, 1, 102, 6, 130, 1, 131, 3, 
/* out0187_had-eta7-phi9*/	3, 63, 4, 102, 2, 130, 3, 
/* out0188_had-eta8-phi9*/	3, 62, 1, 63, 4, 130, 3, 
/* out0189_had-eta9-phi9*/	3, 62, 4, 129, 3, 130, 1, 
/* out0190_had-eta10-phi9*/	3, 15, 1, 62, 3, 129, 5, 
/* out0191_had-eta11-phi9*/	1, 15, 3, 
/* out0192_had-eta12-phi9*/	2, 14, 1, 15, 2, 
/* out0193_had-eta13-phi9*/	1, 14, 2, 
/* out0194_had-eta14-phi9*/	1, 14, 2, 
/* out0195_had-eta15-phi9*/	1, 14, 1, 
/* out0196_had-eta16-phi9*/	1, 18, 1, 
/* out0197_had-eta17-phi9*/	1, 18, 1, 
/* out0198_had-eta18-phi9*/	1, 18, 1, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 133, 4, 
/* out0202_had-eta2-phi10*/	3, 106, 1, 107, 4, 133, 4, 
/* out0203_had-eta3-phi10*/	4, 105, 5, 106, 3, 107, 7, 132, 5, 
/* out0204_had-eta4-phi10*/	5, 65, 2, 103, 1, 105, 8, 131, 1, 132, 3, 
/* out0205_had-eta5-phi10*/	4, 64, 2, 65, 3, 103, 4, 131, 4, 
/* out0206_had-eta6-phi10*/	3, 64, 7, 130, 1, 131, 3, 
/* out0207_had-eta7-phi10*/	3, 63, 4, 64, 2, 130, 3, 
/* out0208_had-eta8-phi10*/	3, 63, 4, 74, 1, 130, 3, 
/* out0209_had-eta9-phi10*/	3, 74, 4, 129, 3, 130, 1, 
/* out0210_had-eta10-phi10*/	3, 15, 2, 74, 2, 129, 5, 
/* out0211_had-eta11-phi10*/	1, 15, 3, 
/* out0212_had-eta12-phi10*/	1, 15, 2, 
/* out0213_had-eta13-phi10*/	2, 14, 1, 19, 1, 
/* out0214_had-eta14-phi10*/	1, 14, 1, 
/* out0215_had-eta15-phi10*/	2, 14, 1, 18, 1, 
/* out0216_had-eta16-phi10*/	1, 18, 1, 
/* out0217_had-eta17-phi10*/	1, 18, 1, 
/* out0218_had-eta18-phi10*/	1, 18, 1, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 138, 4, 
/* out0222_had-eta2-phi11*/	3, 67, 5, 107, 2, 138, 4, 
/* out0223_had-eta3-phi11*/	4, 66, 8, 67, 5, 107, 3, 137, 5, 
/* out0224_had-eta4-phi11*/	5, 65, 5, 66, 6, 77, 1, 136, 1, 137, 3, 
/* out0225_had-eta5-phi11*/	4, 64, 1, 65, 6, 76, 2, 136, 4, 
/* out0226_had-eta6-phi11*/	5, 64, 3, 75, 1, 76, 4, 135, 1, 136, 3, 
/* out0227_had-eta7-phi11*/	2, 75, 6, 135, 3, 
/* out0228_had-eta8-phi11*/	3, 74, 2, 75, 3, 135, 3, 
/* out0229_had-eta9-phi11*/	3, 74, 4, 134, 3, 135, 1, 
/* out0230_had-eta10-phi11*/	3, 20, 1, 74, 2, 134, 5, 
/* out0231_had-eta11-phi11*/	2, 15, 2, 20, 1, 
/* out0232_had-eta12-phi11*/	2, 15, 1, 19, 1, 
/* out0233_had-eta13-phi11*/	1, 19, 2, 
/* out0234_had-eta14-phi11*/	1, 19, 2, 
/* out0235_had-eta15-phi11*/	1, 18, 1, 
/* out0236_had-eta16-phi11*/	1, 18, 1, 
/* out0237_had-eta17-phi11*/	1, 18, 1, 
/* out0238_had-eta18-phi11*/	1, 18, 1, 
/* out0239_had-eta19-phi11*/	1, 18, 1, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 138, 4, 
/* out0242_had-eta2-phi12*/	2, 67, 2, 138, 4, 
/* out0243_had-eta3-phi12*/	4, 66, 1, 67, 4, 78, 9, 137, 5, 
/* out0244_had-eta4-phi12*/	5, 66, 1, 77, 9, 78, 1, 136, 1, 137, 3, 
/* out0245_had-eta5-phi12*/	4, 76, 4, 77, 4, 86, 1, 136, 4, 
/* out0246_had-eta6-phi12*/	4, 76, 6, 85, 1, 135, 1, 136, 3, 
/* out0247_had-eta7-phi12*/	3, 75, 4, 85, 2, 135, 3, 
/* out0248_had-eta8-phi12*/	3, 75, 2, 84, 3, 135, 3, 
/* out0249_had-eta9-phi12*/	4, 74, 1, 84, 3, 134, 3, 135, 1, 
/* out0250_had-eta10-phi12*/	2, 20, 3, 134, 5, 
/* out0251_had-eta11-phi12*/	1, 20, 3, 
/* out0252_had-eta12-phi12*/	2, 19, 1, 20, 1, 
/* out0253_had-eta13-phi12*/	1, 19, 2, 
/* out0254_had-eta14-phi12*/	1, 19, 2, 
/* out0255_had-eta15-phi12*/	1, 19, 1, 
/* out0256_had-eta16-phi12*/	1, 18, 1, 
/* out0257_had-eta17-phi12*/	1, 18, 1, 
/* out0258_had-eta18-phi12*/	1, 18, 1, 
/* out0259_had-eta19-phi12*/	1, 4, 1, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 143, 4, 
/* out0262_had-eta2-phi13*/	1, 143, 4, 
/* out0263_had-eta3-phi13*/	4, 78, 5, 87, 2, 88, 9, 142, 5, 
/* out0264_had-eta4-phi13*/	5, 77, 2, 78, 1, 87, 8, 141, 1, 142, 3, 
/* out0265_had-eta5-phi13*/	2, 86, 8, 141, 4, 
/* out0266_had-eta6-phi13*/	4, 85, 4, 86, 3, 140, 1, 141, 3, 
/* out0267_had-eta7-phi13*/	2, 85, 6, 140, 3, 
/* out0268_had-eta8-phi13*/	2, 84, 5, 140, 3, 
/* out0269_had-eta9-phi13*/	3, 84, 4, 139, 3, 140, 1, 
/* out0270_had-eta10-phi13*/	2, 20, 3, 139, 5, 
/* out0271_had-eta11-phi13*/	1, 20, 3, 
/* out0272_had-eta12-phi13*/	3, 7, 1, 19, 1, 20, 1, 
/* out0273_had-eta13-phi13*/	1, 19, 2, 
/* out0274_had-eta14-phi13*/	1, 19, 1, 
/* out0275_had-eta15-phi13*/	1, 6, 1, 
/* out0276_had-eta16-phi13*/	1, 6, 1, 
/* out0277_had-eta17-phi13*/	1, 18, 1, 
/* out0278_had-eta18-phi13*/	1, 4, 2, 
/* out0279_had-eta19-phi13*/	1, 4, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 143, 4, 
/* out0282_had-eta2-phi14*/	1, 143, 4, 
/* out0283_had-eta3-phi14*/	3, 87, 1, 88, 7, 142, 5, 
/* out0284_had-eta4-phi14*/	4, 31, 4, 87, 5, 141, 1, 142, 3, 
/* out0285_had-eta5-phi14*/	4, 30, 1, 31, 4, 86, 3, 141, 4, 
/* out0286_had-eta6-phi14*/	5, 30, 6, 85, 1, 86, 1, 140, 1, 141, 3, 
/* out0287_had-eta7-phi14*/	4, 29, 3, 30, 1, 85, 2, 140, 3, 
/* out0288_had-eta8-phi14*/	2, 29, 5, 140, 3, 
/* out0289_had-eta9-phi14*/	4, 28, 3, 84, 1, 139, 3, 140, 1, 
/* out0290_had-eta10-phi14*/	2, 28, 3, 139, 5, 
/* out0291_had-eta11-phi14*/	2, 7, 2, 28, 1, 
/* out0292_had-eta12-phi14*/	1, 7, 2, 
/* out0293_had-eta13-phi14*/	1, 7, 2, 
/* out0294_had-eta14-phi14*/	1, 6, 2, 
/* out0295_had-eta15-phi14*/	1, 6, 1, 
/* out0296_had-eta16-phi14*/	1, 6, 1, 
/* out0297_had-eta17-phi14*/	1, 6, 1, 
/* out0298_had-eta18-phi14*/	1, 4, 2, 
/* out0299_had-eta19-phi14*/	1, 4, 2, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 148, 4, 
/* out0302_had-eta2-phi15*/	1, 148, 4, 
/* out0303_had-eta3-phi15*/	3, 40, 1, 41, 7, 147, 5, 
/* out0304_had-eta4-phi15*/	4, 31, 4, 40, 5, 146, 1, 147, 3, 
/* out0305_had-eta5-phi15*/	4, 30, 1, 31, 4, 39, 3, 146, 4, 
/* out0306_had-eta6-phi15*/	5, 30, 6, 38, 1, 39, 1, 145, 1, 146, 3, 
/* out0307_had-eta7-phi15*/	4, 29, 3, 30, 1, 38, 2, 145, 3, 
/* out0308_had-eta8-phi15*/	2, 29, 5, 145, 3, 
/* out0309_had-eta9-phi15*/	4, 28, 3, 37, 1, 144, 3, 145, 1, 
/* out0310_had-eta10-phi15*/	2, 28, 4, 144, 5, 
/* out0311_had-eta11-phi15*/	2, 7, 2, 28, 1, 
/* out0312_had-eta12-phi15*/	1, 7, 3, 
/* out0313_had-eta13-phi15*/	1, 7, 2, 
/* out0314_had-eta14-phi15*/	1, 6, 2, 
/* out0315_had-eta15-phi15*/	1, 6, 1, 
/* out0316_had-eta16-phi15*/	1, 6, 1, 
/* out0317_had-eta17-phi15*/	1, 6, 1, 
/* out0318_had-eta18-phi15*/	1, 4, 2, 
/* out0319_had-eta19-phi15*/	1, 4, 2, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 148, 4, 
/* out0322_had-eta2-phi16*/	1, 148, 4, 
/* out0323_had-eta3-phi16*/	4, 40, 2, 41, 9, 51, 5, 147, 5, 
/* out0324_had-eta4-phi16*/	5, 40, 8, 50, 2, 51, 1, 146, 1, 147, 3, 
/* out0325_had-eta5-phi16*/	2, 39, 8, 146, 4, 
/* out0326_had-eta6-phi16*/	4, 38, 4, 39, 3, 145, 1, 146, 3, 
/* out0327_had-eta7-phi16*/	2, 38, 6, 145, 3, 
/* out0328_had-eta8-phi16*/	2, 37, 5, 145, 3, 
/* out0329_had-eta9-phi16*/	3, 37, 4, 144, 3, 145, 1, 
/* out0330_had-eta10-phi16*/	3, 13, 3, 28, 1, 144, 5, 
/* out0331_had-eta11-phi16*/	1, 13, 3, 
/* out0332_had-eta12-phi16*/	3, 7, 1, 11, 1, 13, 1, 
/* out0333_had-eta13-phi16*/	2, 7, 1, 11, 2, 
/* out0334_had-eta14-phi16*/	2, 6, 1, 11, 1, 
/* out0335_had-eta15-phi16*/	1, 6, 1, 
/* out0336_had-eta16-phi16*/	1, 6, 1, 
/* out0337_had-eta17-phi16*/	2, 5, 1, 6, 1, 
/* out0338_had-eta18-phi16*/	1, 4, 2, 
/* out0339_had-eta19-phi16*/	1, 4, 1, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 153, 4, 
/* out0342_had-eta2-phi17*/	2, 61, 2, 153, 4, 
/* out0343_had-eta3-phi17*/	4, 51, 9, 60, 2, 61, 4, 152, 5, 
/* out0344_had-eta4-phi17*/	5, 50, 9, 51, 1, 60, 1, 151, 1, 152, 3, 
/* out0345_had-eta5-phi17*/	4, 39, 1, 49, 4, 50, 4, 151, 4, 
/* out0346_had-eta6-phi17*/	4, 38, 1, 49, 6, 150, 1, 151, 3, 
/* out0347_had-eta7-phi17*/	3, 38, 2, 48, 4, 150, 3, 
/* out0348_had-eta8-phi17*/	3, 37, 3, 48, 2, 150, 3, 
/* out0349_had-eta9-phi17*/	4, 37, 3, 47, 1, 149, 3, 150, 1, 
/* out0350_had-eta10-phi17*/	2, 13, 3, 149, 5, 
/* out0351_had-eta11-phi17*/	1, 13, 3, 
/* out0352_had-eta12-phi17*/	2, 11, 1, 13, 1, 
/* out0353_had-eta13-phi17*/	1, 11, 2, 
/* out0354_had-eta14-phi17*/	1, 11, 2, 
/* out0355_had-eta15-phi17*/	1, 11, 1, 
/* out0356_had-eta16-phi17*/	1, 5, 1, 
/* out0357_had-eta17-phi17*/	1, 5, 1, 
/* out0358_had-eta18-phi17*/	1, 5, 1, 
/* out0359_had-eta19-phi17*/	1, 4, 1, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 153, 4, 
/* out0362_had-eta2-phi18*/	3, 61, 5, 101, 2, 153, 4, 
/* out0363_had-eta3-phi18*/	4, 60, 8, 61, 5, 101, 3, 152, 5, 
/* out0364_had-eta4-phi18*/	5, 50, 1, 59, 5, 60, 5, 151, 1, 152, 3, 
/* out0365_had-eta5-phi18*/	4, 49, 2, 58, 1, 59, 6, 151, 4, 
/* out0366_had-eta6-phi18*/	5, 48, 1, 49, 4, 58, 3, 150, 1, 151, 3, 
/* out0367_had-eta7-phi18*/	2, 48, 6, 150, 3, 
/* out0368_had-eta8-phi18*/	3, 47, 2, 48, 3, 150, 3, 
/* out0369_had-eta9-phi18*/	3, 47, 4, 149, 3, 150, 1, 
/* out0370_had-eta10-phi18*/	3, 13, 1, 47, 2, 149, 5, 
/* out0371_had-eta11-phi18*/	2, 12, 2, 13, 1, 
/* out0372_had-eta12-phi18*/	2, 11, 1, 12, 1, 
/* out0373_had-eta13-phi18*/	1, 11, 2, 
/* out0374_had-eta14-phi18*/	1, 11, 2, 
/* out0375_had-eta15-phi18*/	1, 5, 1, 
/* out0376_had-eta16-phi18*/	1, 5, 1, 
/* out0377_had-eta17-phi18*/	1, 5, 1, 
/* out0378_had-eta18-phi18*/	1, 5, 1, 
/* out0379_had-eta19-phi18*/	1, 5, 1, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 158, 4, 
/* out0382_had-eta2-phi19*/	3, 100, 1, 101, 4, 158, 4, 
/* out0383_had-eta3-phi19*/	4, 99, 5, 100, 3, 101, 7, 157, 5, 
/* out0384_had-eta4-phi19*/	5, 59, 2, 98, 1, 99, 8, 156, 1, 157, 3, 
/* out0385_had-eta5-phi19*/	4, 58, 2, 59, 3, 98, 4, 156, 4, 
/* out0386_had-eta6-phi19*/	3, 58, 7, 155, 1, 156, 3, 
/* out0387_had-eta7-phi19*/	3, 57, 4, 58, 2, 155, 3, 
/* out0388_had-eta8-phi19*/	3, 47, 1, 57, 4, 155, 3, 
/* out0389_had-eta9-phi19*/	3, 47, 4, 154, 3, 155, 1, 
/* out0390_had-eta10-phi19*/	3, 12, 2, 47, 2, 154, 5, 
/* out0391_had-eta11-phi19*/	1, 12, 3, 
/* out0392_had-eta12-phi19*/	1, 12, 2, 
/* out0393_had-eta13-phi19*/	2, 11, 1, 16, 1, 
/* out0394_had-eta14-phi19*/	1, 16, 1, 
/* out0395_had-eta15-phi19*/	1, 5, 1, 
/* out0396_had-eta16-phi19*/	1, 5, 1, 
/* out0397_had-eta17-phi19*/	1, 5, 1, 
/* out0398_had-eta18-phi19*/	1, 5, 1, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 158, 4, 
/* out0402_had-eta2-phi20*/	1, 158, 4, 
/* out0403_had-eta3-phi20*/	4, 99, 1, 100, 12, 112, 3, 157, 5, 
/* out0404_had-eta4-phi20*/	5, 98, 3, 99, 2, 112, 5, 156, 1, 157, 3, 
/* out0405_had-eta5-phi20*/	2, 98, 8, 156, 4, 
/* out0406_had-eta6-phi20*/	4, 58, 1, 108, 6, 155, 1, 156, 3, 
/* out0407_had-eta7-phi20*/	3, 57, 4, 108, 1, 155, 3, 
/* out0408_had-eta8-phi20*/	3, 57, 4, 68, 1, 155, 3, 
/* out0409_had-eta9-phi20*/	3, 68, 4, 154, 3, 155, 1, 
/* out0410_had-eta10-phi20*/	3, 12, 1, 68, 3, 154, 5, 
/* out0411_had-eta11-phi20*/	1, 12, 3, 
/* out0412_had-eta12-phi20*/	1, 12, 2, 
/* out0413_had-eta13-phi20*/	1, 16, 2, 
/* out0414_had-eta14-phi20*/	1, 16, 2, 
/* out0415_had-eta15-phi20*/	1, 16, 1, 
/* out0416_had-eta16-phi20*/	1, 5, 1, 
/* out0417_had-eta17-phi20*/	1, 5, 1, 
/* out0418_had-eta18-phi20*/	1, 5, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 163, 4, 
/* out0422_had-eta2-phi21*/	1, 163, 4, 
/* out0423_had-eta3-phi21*/	4, 110, 1, 112, 3, 113, 12, 162, 5, 
/* out0424_had-eta4-phi21*/	5, 109, 3, 110, 2, 112, 5, 161, 1, 162, 3, 
/* out0425_had-eta5-phi21*/	3, 108, 1, 109, 8, 161, 4, 
/* out0426_had-eta6-phi21*/	4, 70, 1, 108, 6, 160, 1, 161, 3, 
/* out0427_had-eta7-phi21*/	3, 69, 4, 108, 2, 160, 3, 
/* out0428_had-eta8-phi21*/	3, 68, 1, 69, 4, 160, 3, 
/* out0429_had-eta9-phi21*/	3, 68, 4, 159, 3, 160, 1, 
/* out0430_had-eta10-phi21*/	3, 17, 1, 68, 3, 159, 5, 
/* out0431_had-eta11-phi21*/	1, 17, 3, 
/* out0432_had-eta12-phi21*/	2, 16, 1, 17, 2, 
/* out0433_had-eta13-phi21*/	1, 16, 2, 
/* out0434_had-eta14-phi21*/	1, 16, 2, 
/* out0435_had-eta15-phi21*/	1, 16, 1, 
/* out0436_had-eta16-phi21*/	1, 21, 1, 
/* out0437_had-eta17-phi21*/	1, 21, 1, 
/* out0438_had-eta18-phi21*/	1, 21, 1, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 163, 4, 
/* out0442_had-eta2-phi22*/	3, 111, 4, 113, 1, 163, 4, 
/* out0443_had-eta3-phi22*/	4, 110, 5, 111, 7, 113, 3, 162, 5, 
/* out0444_had-eta4-phi22*/	5, 71, 2, 109, 1, 110, 8, 161, 1, 162, 3, 
/* out0445_had-eta5-phi22*/	4, 70, 2, 71, 3, 109, 4, 161, 4, 
/* out0446_had-eta6-phi22*/	3, 70, 7, 160, 1, 161, 3, 
/* out0447_had-eta7-phi22*/	3, 69, 4, 70, 2, 160, 3, 
/* out0448_had-eta8-phi22*/	3, 69, 4, 79, 1, 160, 3, 
/* out0449_had-eta9-phi22*/	3, 79, 4, 159, 3, 160, 1, 
/* out0450_had-eta10-phi22*/	3, 17, 2, 79, 2, 159, 5, 
/* out0451_had-eta11-phi22*/	1, 17, 3, 
/* out0452_had-eta12-phi22*/	1, 17, 2, 
/* out0453_had-eta13-phi22*/	2, 16, 1, 22, 1, 
/* out0454_had-eta14-phi22*/	1, 16, 1, 
/* out0455_had-eta15-phi22*/	2, 16, 1, 21, 1, 
/* out0456_had-eta16-phi22*/	1, 21, 1, 
/* out0457_had-eta17-phi22*/	1, 21, 1, 
/* out0458_had-eta18-phi22*/	1, 21, 1, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 168, 4, 
/* out0462_had-eta2-phi23*/	3, 73, 5, 111, 2, 168, 4, 
/* out0463_had-eta3-phi23*/	4, 72, 8, 73, 5, 111, 3, 167, 5, 
/* out0464_had-eta4-phi23*/	5, 71, 5, 72, 5, 82, 1, 166, 1, 167, 3, 
/* out0465_had-eta5-phi23*/	4, 70, 1, 71, 6, 81, 2, 166, 4, 
/* out0466_had-eta6-phi23*/	5, 70, 3, 80, 1, 81, 4, 165, 1, 166, 3, 
/* out0467_had-eta7-phi23*/	2, 80, 6, 165, 3, 
/* out0468_had-eta8-phi23*/	3, 79, 2, 80, 3, 165, 3, 
/* out0469_had-eta9-phi23*/	3, 79, 4, 164, 3, 165, 1, 
/* out0470_had-eta10-phi23*/	3, 23, 1, 79, 2, 164, 5, 
/* out0471_had-eta11-phi23*/	2, 17, 2, 23, 1, 
/* out0472_had-eta12-phi23*/	2, 17, 1, 22, 1, 
/* out0473_had-eta13-phi23*/	1, 22, 2, 
/* out0474_had-eta14-phi23*/	1, 22, 2, 
/* out0475_had-eta15-phi23*/	1, 21, 1, 
/* out0476_had-eta16-phi23*/	1, 21, 1, 
/* out0477_had-eta17-phi23*/	1, 21, 1, 
/* out0478_had-eta18-phi23*/	1, 21, 1, 
/* out0479_had-eta19-phi23*/	1, 21, 1, 
/* out0480_had-eta0-phi24*/	0, 
/* out0481_had-eta1-phi24*/	1, 168, 4, 
/* out0482_had-eta2-phi24*/	2, 73, 2, 168, 4, 
/* out0483_had-eta3-phi24*/	4, 72, 2, 73, 4, 83, 9, 167, 5, 
/* out0484_had-eta4-phi24*/	5, 72, 1, 82, 9, 83, 1, 166, 1, 167, 3, 
/* out0485_had-eta5-phi24*/	4, 81, 4, 82, 4, 91, 1, 166, 4, 
/* out0486_had-eta6-phi24*/	4, 81, 6, 90, 1, 165, 1, 166, 3, 
/* out0487_had-eta7-phi24*/	3, 80, 4, 90, 2, 165, 3, 
/* out0488_had-eta8-phi24*/	3, 80, 2, 89, 3, 165, 3, 
/* out0489_had-eta9-phi24*/	4, 79, 1, 89, 3, 164, 3, 165, 1, 
/* out0490_had-eta10-phi24*/	2, 23, 3, 164, 5, 
/* out0491_had-eta11-phi24*/	1, 23, 3, 
/* out0492_had-eta12-phi24*/	2, 22, 1, 23, 1, 
/* out0493_had-eta13-phi24*/	1, 22, 2, 
/* out0494_had-eta14-phi24*/	1, 22, 2, 
/* out0495_had-eta15-phi24*/	1, 22, 1, 
/* out0496_had-eta16-phi24*/	1, 21, 1, 
/* out0497_had-eta17-phi24*/	1, 21, 1, 
/* out0498_had-eta18-phi24*/	1, 21, 1, 
/* out0499_had-eta19-phi24*/	0, 
/* out0500_had-eta0-phi25*/	0, 
/* out0501_had-eta1-phi25*/	1, 173, 4, 
/* out0502_had-eta2-phi25*/	1, 173, 4, 
/* out0503_had-eta3-phi25*/	4, 83, 5, 92, 2, 93, 9, 172, 5, 
/* out0504_had-eta4-phi25*/	5, 82, 2, 83, 1, 92, 8, 171, 1, 172, 3, 
/* out0505_had-eta5-phi25*/	2, 91, 8, 171, 4, 
/* out0506_had-eta6-phi25*/	4, 90, 4, 91, 3, 170, 1, 171, 3, 
/* out0507_had-eta7-phi25*/	2, 90, 6, 170, 3, 
/* out0508_had-eta8-phi25*/	2, 89, 5, 170, 3, 
/* out0509_had-eta9-phi25*/	3, 89, 4, 169, 3, 170, 1, 
/* out0510_had-eta10-phi25*/	2, 23, 3, 169, 5, 
/* out0511_had-eta11-phi25*/	1, 23, 3, 
/* out0512_had-eta12-phi25*/	2, 22, 1, 23, 1, 
/* out0513_had-eta13-phi25*/	1, 22, 2, 
/* out0514_had-eta14-phi25*/	1, 22, 1, 
/* out0515_had-eta15-phi25*/	0, 
/* out0516_had-eta16-phi25*/	0, 
/* out0517_had-eta17-phi25*/	1, 21, 1, 
/* out0518_had-eta18-phi25*/	0, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	0, 
/* out0521_had-eta1-phi26*/	1, 173, 4, 
/* out0522_had-eta2-phi26*/	1, 173, 4, 
/* out0523_had-eta3-phi26*/	3, 92, 1, 93, 7, 172, 5, 
/* out0524_had-eta4-phi26*/	3, 92, 5, 171, 1, 172, 3, 
/* out0525_had-eta5-phi26*/	2, 91, 3, 171, 4, 
/* out0526_had-eta6-phi26*/	4, 90, 1, 91, 1, 170, 1, 171, 3, 
/* out0527_had-eta7-phi26*/	2, 90, 2, 170, 3, 
/* out0528_had-eta8-phi26*/	1, 170, 3, 
/* out0529_had-eta9-phi26*/	3, 89, 1, 169, 3, 170, 1, 
/* out0530_had-eta10-phi26*/	1, 169, 5, 
/* out0531_had-eta11-phi26*/	0, 
/* out0532_had-eta12-phi26*/	0, 
/* out0533_had-eta13-phi26*/	0, 
/* out0534_had-eta14-phi26*/	0, 
/* out0535_had-eta15-phi26*/	0, 
/* out0536_had-eta16-phi26*/	0, 
/* out0537_had-eta17-phi26*/	0, 
/* out0538_had-eta18-phi26*/	0, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	0, 
/* out0550_had-eta10-phi27*/	0, 
/* out0551_had-eta11-phi27*/	0, 
/* out0552_had-eta12-phi27*/	0, 
/* out0553_had-eta13-phi27*/	0, 
/* out0554_had-eta14-phi27*/	0, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	0, 
/* out0557_had-eta17-phi27*/	0, 
/* out0558_had-eta18-phi27*/	0, 
/* out0559_had-eta19-phi27*/	0, 
};