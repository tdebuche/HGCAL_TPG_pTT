parameter integer matrixH [0:6137] = {
/* num inputs = 174(in0-in173) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1859 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	1, 0, 6, 4, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	1, 24, 2, 1, 
/* out0030_had-eta10-phi1*/	1, 24, 1, 1, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	2, 3, 5, 6, 3, 11, 7, 
/* out0033_had-eta13-phi1*/	2, 3, 4, 2, 3, 5, 3, 
/* out0034_had-eta14-phi1*/	2, 1, 8, 3, 1, 11, 1, 
/* out0035_had-eta15-phi1*/	2, 1, 5, 4, 1, 11, 11, 
/* out0036_had-eta16-phi1*/	2, 1, 4, 2, 1, 5, 9, 
/* out0037_had-eta17-phi1*/	2, 0, 3, 1, 1, 4, 5, 
/* out0038_had-eta18-phi1*/	1, 0, 3, 7, 
/* out0039_had-eta19-phi1*/	1, 0, 6, 11, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	1, 27, 2, 11, 
/* out0045_had-eta5-phi2*/	3, 26, 2, 4, 27, 1, 12, 27, 2, 1, 
/* out0046_had-eta6-phi2*/	2, 26, 1, 9, 26, 2, 8, 
/* out0047_had-eta7-phi2*/	2, 25, 2, 10, 26, 1, 3, 
/* out0048_had-eta8-phi2*/	2, 25, 1, 11, 25, 2, 2, 
/* out0049_had-eta9-phi2*/	2, 24, 2, 9, 25, 1, 1, 
/* out0050_had-eta10-phi2*/	2, 24, 1, 9, 24, 2, 2, 
/* out0051_had-eta11-phi2*/	4, 3, 8, 16, 3, 9, 4, 3, 11, 1, 24, 1, 2, 
/* out0052_had-eta12-phi2*/	4, 3, 5, 3, 3, 6, 7, 3, 10, 11, 3, 11, 8, 
/* out0053_had-eta13-phi2*/	4, 3, 4, 11, 3, 5, 4, 3, 6, 5, 3, 7, 3, 
/* out0054_had-eta14-phi2*/	4, 1, 8, 13, 1, 9, 4, 1, 11, 1, 3, 4, 3, 
/* out0055_had-eta15-phi2*/	3, 1, 6, 2, 1, 10, 11, 1, 11, 3, 
/* out0056_had-eta16-phi2*/	4, 1, 4, 1, 1, 5, 3, 1, 6, 9, 1, 7, 1, 
/* out0057_had-eta17-phi2*/	3, 0, 3, 1, 1, 4, 8, 1, 7, 3, 
/* out0058_had-eta18-phi2*/	2, 0, 3, 7, 0, 4, 3, 
/* out0059_had-eta19-phi2*/	2, 0, 5, 10, 0, 6, 1, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 118, 0, 4, 
/* out0062_had-eta2-phi3*/	1, 118, 0, 4, 
/* out0063_had-eta3-phi3*/	3, 35, 2, 3, 36, 1, 10, 117, 0, 5, 
/* out0064_had-eta4-phi3*/	6, 27, 0, 8, 27, 2, 4, 35, 1, 8, 35, 2, 6, 116, 0, 1, 117, 0, 3, 
/* out0065_had-eta5-phi3*/	7, 26, 0, 1, 26, 2, 2, 27, 0, 8, 27, 1, 4, 34, 1, 3, 34, 2, 7, 116, 0, 4, 
/* out0066_had-eta6-phi3*/	7, 26, 0, 14, 26, 1, 2, 26, 2, 2, 33, 2, 2, 34, 1, 2, 115, 0, 1, 116, 0, 3, 
/* out0067_had-eta7-phi3*/	7, 25, 0, 6, 25, 2, 4, 26, 0, 1, 26, 1, 2, 33, 1, 3, 33, 2, 2, 115, 0, 3, 
/* out0068_had-eta8-phi3*/	4, 25, 0, 10, 25, 1, 3, 32, 2, 2, 115, 0, 3, 
/* out0069_had-eta9-phi3*/	6, 24, 0, 5, 24, 2, 4, 25, 1, 1, 32, 1, 2, 114, 0, 3, 115, 0, 1, 
/* out0070_had-eta10-phi3*/	3, 24, 0, 8, 24, 1, 2, 114, 0, 5, 
/* out0071_had-eta11-phi3*/	7, 3, 3, 8, 3, 9, 12, 3, 10, 1, 9, 1, 1, 9, 2, 1, 24, 0, 1, 24, 1, 2, 
/* out0072_had-eta12-phi3*/	6, 3, 0, 1, 3, 1, 2, 3, 2, 14, 3, 3, 6, 3, 6, 1, 3, 10, 4, 
/* out0073_had-eta13-phi3*/	4, 3, 1, 9, 3, 2, 2, 3, 6, 3, 3, 7, 10, 
/* out0074_had-eta14-phi3*/	4, 1, 3, 4, 1, 9, 12, 1, 10, 1, 3, 7, 3, 
/* out0075_had-eta15-phi3*/	3, 1, 2, 10, 1, 3, 3, 1, 10, 4, 
/* out0076_had-eta16-phi3*/	4, 1, 1, 3, 1, 2, 6, 1, 6, 5, 1, 7, 1, 
/* out0077_had-eta17-phi3*/	3, 0, 4, 1, 1, 1, 1, 1, 7, 10, 
/* out0078_had-eta18-phi3*/	2, 0, 2, 1, 0, 4, 10, 
/* out0079_had-eta19-phi3*/	4, 0, 1, 14, 0, 2, 1, 0, 4, 1, 0, 5, 6, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 118, 0, 4, 
/* out0082_had-eta2-phi4*/	1, 118, 0, 4, 
/* out0083_had-eta3-phi4*/	7, 35, 0, 2, 35, 2, 4, 36, 0, 16, 36, 1, 6, 46, 1, 5, 46, 2, 9, 117, 0, 5, 
/* out0084_had-eta4-phi4*/	9, 34, 2, 1, 35, 0, 14, 35, 1, 8, 35, 2, 3, 45, 1, 1, 45, 2, 4, 46, 1, 1, 116, 0, 1, 117, 0, 3, 
/* out0085_had-eta5-phi4*/	5, 34, 0, 13, 34, 1, 4, 34, 2, 8, 45, 1, 1, 116, 0, 4, 
/* out0086_had-eta6-phi4*/	7, 33, 0, 3, 33, 2, 10, 34, 0, 1, 34, 1, 7, 44, 2, 1, 115, 0, 1, 116, 0, 3, 
/* out0087_had-eta7-phi4*/	4, 33, 0, 4, 33, 1, 12, 33, 2, 2, 115, 0, 3, 
/* out0088_had-eta8-phi4*/	4, 32, 0, 1, 32, 2, 13, 33, 1, 1, 115, 0, 3, 
/* out0089_had-eta9-phi4*/	3, 32, 1, 11, 114, 0, 3, 115, 0, 1, 
/* out0090_had-eta10-phi4*/	3, 9, 2, 9, 24, 0, 2, 114, 0, 5, 
/* out0091_had-eta11-phi4*/	3, 3, 3, 1, 9, 1, 6, 9, 2, 2, 
/* out0092_had-eta12-phi4*/	4, 3, 0, 13, 3, 3, 1, 8, 8, 6, 9, 1, 2, 
/* out0093_had-eta13-phi4*/	4, 3, 0, 2, 3, 1, 5, 8, 8, 4, 8, 11, 14, 
/* out0094_had-eta14-phi4*/	4, 1, 3, 5, 8, 4, 1, 8, 5, 13, 8, 11, 1, 
/* out0095_had-eta15-phi4*/	3, 1, 0, 11, 1, 3, 4, 8, 4, 2, 
/* out0096_had-eta16-phi4*/	4, 1, 0, 4, 1, 1, 8, 2, 8, 1, 2, 11, 1, 
/* out0097_had-eta17-phi4*/	4, 1, 1, 4, 1, 7, 1, 2, 5, 1, 2, 11, 4, 
/* out0098_had-eta18-phi4*/	3, 0, 2, 8, 0, 4, 1, 2, 5, 2, 
/* out0099_had-eta19-phi4*/	3, 0, 0, 1, 0, 1, 2, 0, 2, 6, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 123, 0, 4, 
/* out0102_had-eta2-phi5*/	2, 56, 1, 2, 123, 0, 4, 
/* out0103_had-eta3-phi5*/	6, 46, 0, 16, 46, 1, 6, 46, 2, 7, 55, 2, 4, 56, 1, 7, 122, 0, 5, 
/* out0104_had-eta4-phi5*/	8, 45, 0, 11, 45, 1, 3, 45, 2, 12, 46, 1, 4, 55, 1, 2, 55, 2, 1, 121, 0, 1, 122, 0, 3, 
/* out0105_had-eta5-phi5*/	6, 34, 0, 2, 44, 0, 1, 44, 2, 11, 45, 0, 2, 45, 1, 11, 121, 0, 4, 
/* out0106_had-eta6-phi5*/	7, 33, 0, 3, 43, 2, 1, 44, 0, 1, 44, 1, 13, 44, 2, 4, 120, 0, 1, 121, 0, 3, 
/* out0107_had-eta7-phi5*/	4, 33, 0, 6, 43, 1, 2, 43, 2, 10, 120, 0, 3, 
/* out0108_had-eta8-phi5*/	4, 32, 0, 9, 32, 2, 1, 43, 1, 5, 120, 0, 3, 
/* out0109_had-eta9-phi5*/	6, 32, 0, 6, 32, 1, 3, 42, 1, 1, 42, 2, 3, 119, 0, 3, 120, 0, 1, 
/* out0110_had-eta10-phi5*/	3, 9, 0, 6, 9, 2, 4, 119, 0, 5, 
/* out0111_had-eta11-phi5*/	2, 9, 0, 4, 9, 1, 4, 
/* out0112_had-eta12-phi5*/	3, 8, 8, 5, 8, 9, 12, 9, 1, 3, 
/* out0113_had-eta13-phi5*/	6, 8, 2, 3, 8, 6, 2, 8, 8, 1, 8, 9, 2, 8, 10, 16, 8, 11, 1, 
/* out0114_had-eta14-phi5*/	4, 8, 4, 3, 8, 5, 3, 8, 6, 11, 8, 7, 3, 
/* out0115_had-eta15-phi5*/	4, 1, 0, 1, 2, 8, 6, 8, 4, 10, 8, 7, 1, 
/* out0116_had-eta16-phi5*/	3, 2, 8, 8, 2, 10, 1, 2, 11, 5, 
/* out0117_had-eta17-phi5*/	4, 2, 5, 3, 2, 6, 1, 2, 10, 2, 2, 11, 6, 
/* out0118_had-eta18-phi5*/	2, 2, 4, 2, 2, 5, 8, 
/* out0119_had-eta19-phi5*/	2, 0, 0, 15, 2, 4, 2, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 123, 0, 4, 
/* out0122_had-eta2-phi6*/	4, 56, 0, 12, 56, 1, 1, 96, 2, 7, 123, 0, 4, 
/* out0123_had-eta3-phi6*/	8, 55, 0, 12, 55, 1, 1, 55, 2, 11, 56, 0, 4, 56, 1, 6, 96, 1, 5, 96, 2, 4, 122, 0, 5, 
/* out0124_had-eta4-phi6*/	7, 45, 0, 3, 54, 0, 2, 54, 2, 11, 55, 0, 3, 55, 1, 13, 121, 0, 1, 122, 0, 3, 
/* out0125_had-eta5-phi6*/	6, 44, 0, 6, 53, 2, 1, 54, 0, 1, 54, 1, 13, 54, 2, 5, 121, 0, 4, 
/* out0126_had-eta6-phi6*/	8, 43, 0, 1, 43, 2, 1, 44, 0, 8, 44, 1, 3, 53, 1, 3, 53, 2, 7, 120, 0, 1, 121, 0, 3, 
/* out0127_had-eta7-phi6*/	5, 43, 0, 11, 43, 1, 2, 43, 2, 4, 53, 1, 1, 120, 0, 3, 
/* out0128_had-eta8-phi6*/	4, 42, 2, 6, 43, 0, 2, 43, 1, 7, 120, 0, 3, 
/* out0129_had-eta9-phi6*/	5, 42, 0, 1, 42, 1, 4, 42, 2, 7, 119, 0, 3, 120, 0, 1, 
/* out0130_had-eta10-phi6*/	4, 9, 0, 3, 10, 8, 5, 42, 1, 7, 119, 0, 5, 
/* out0131_had-eta11-phi6*/	3, 9, 0, 3, 10, 8, 8, 10, 11, 13, 
/* out0132_had-eta12-phi6*/	6, 8, 0, 1, 8, 3, 11, 8, 9, 2, 10, 4, 1, 10, 5, 10, 10, 11, 2, 
/* out0133_had-eta13-phi6*/	4, 8, 0, 6, 8, 1, 3, 8, 2, 10, 8, 3, 5, 
/* out0134_had-eta14-phi6*/	4, 8, 1, 8, 8, 2, 3, 8, 6, 3, 8, 7, 7, 
/* out0135_had-eta15-phi6*/	3, 2, 8, 1, 2, 9, 10, 8, 7, 5, 
/* out0136_had-eta16-phi6*/	3, 2, 2, 1, 2, 9, 4, 2, 10, 9, 
/* out0137_had-eta17-phi6*/	3, 2, 2, 1, 2, 6, 7, 2, 10, 4, 
/* out0138_had-eta18-phi6*/	4, 2, 4, 3, 2, 5, 2, 2, 6, 4, 2, 7, 1, 
/* out0139_had-eta19-phi6*/	1, 2, 4, 7, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 128, 0, 4, 
/* out0142_had-eta2-phi7*/	4, 96, 0, 8, 96, 2, 4, 97, 1, 2, 128, 0, 4, 
/* out0143_had-eta3-phi7*/	9, 55, 0, 1, 95, 0, 5, 95, 2, 10, 96, 0, 8, 96, 1, 11, 96, 2, 1, 97, 0, 1, 97, 1, 7, 127, 0, 5, 
/* out0144_had-eta4-phi7*/	7, 54, 0, 6, 94, 2, 3, 95, 0, 2, 95, 1, 14, 95, 2, 6, 126, 0, 1, 127, 0, 3, 
/* out0145_had-eta5-phi7*/	7, 53, 0, 3, 53, 2, 3, 54, 0, 7, 54, 1, 3, 94, 1, 4, 94, 2, 7, 126, 0, 4, 
/* out0146_had-eta6-phi7*/	5, 53, 0, 10, 53, 1, 7, 53, 2, 5, 125, 0, 1, 126, 0, 3, 
/* out0147_had-eta7-phi7*/	4, 43, 0, 2, 52, 2, 11, 53, 1, 5, 125, 0, 3, 
/* out0148_had-eta8-phi7*/	4, 42, 0, 3, 52, 1, 8, 52, 2, 3, 125, 0, 3, 
/* out0149_had-eta9-phi7*/	5, 42, 0, 11, 42, 1, 1, 62, 2, 1, 124, 0, 3, 125, 0, 1, 
/* out0150_had-eta10-phi7*/	6, 10, 3, 5, 10, 8, 2, 10, 9, 13, 42, 0, 1, 42, 1, 3, 124, 0, 5, 
/* out0151_had-eta11-phi7*/	7, 10, 2, 8, 10, 3, 1, 10, 6, 6, 10, 8, 1, 10, 9, 3, 10, 10, 16, 10, 11, 1, 
/* out0152_had-eta12-phi7*/	4, 10, 4, 11, 10, 5, 6, 10, 6, 9, 10, 7, 3, 
/* out0153_had-eta13-phi7*/	3, 8, 0, 9, 10, 4, 3, 14, 8, 10, 
/* out0154_had-eta14-phi7*/	3, 8, 1, 5, 14, 5, 1, 14, 11, 11, 
/* out0155_had-eta15-phi7*/	3, 2, 3, 9, 2, 9, 2, 14, 5, 5, 
/* out0156_had-eta16-phi7*/	3, 2, 0, 1, 2, 2, 6, 2, 3, 7, 
/* out0157_had-eta17-phi7*/	3, 2, 1, 2, 2, 2, 8, 2, 6, 2, 
/* out0158_had-eta18-phi7*/	2, 2, 6, 2, 2, 7, 8, 
/* out0159_had-eta19-phi7*/	2, 2, 4, 2, 2, 7, 2, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 128, 0, 4, 
/* out0162_had-eta2-phi8*/	1, 128, 0, 4, 
/* out0163_had-eta3-phi8*/	5, 95, 0, 4, 97, 0, 15, 97, 1, 7, 104, 2, 8, 127, 0, 5, 
/* out0164_had-eta4-phi8*/	8, 94, 0, 6, 94, 2, 3, 95, 0, 5, 95, 1, 2, 104, 1, 8, 104, 2, 8, 126, 0, 1, 127, 0, 3, 
/* out0165_had-eta5-phi8*/	5, 94, 0, 10, 94, 1, 11, 94, 2, 3, 102, 2, 2, 126, 0, 4, 
/* out0166_had-eta6-phi8*/	6, 53, 0, 3, 94, 1, 1, 102, 1, 3, 102, 2, 14, 125, 0, 1, 126, 0, 3, 
/* out0167_had-eta7-phi8*/	4, 52, 0, 12, 52, 2, 2, 102, 1, 4, 125, 0, 3, 
/* out0168_had-eta8-phi8*/	4, 52, 0, 4, 52, 1, 8, 62, 2, 2, 125, 0, 3, 
/* out0169_had-eta9-phi8*/	4, 62, 1, 1, 62, 2, 12, 124, 0, 3, 125, 0, 1, 
/* out0170_had-eta10-phi8*/	5, 10, 0, 3, 10, 3, 6, 62, 1, 7, 62, 2, 1, 124, 0, 5, 
/* out0171_had-eta11-phi8*/	4, 10, 0, 13, 10, 1, 9, 10, 2, 8, 10, 3, 4, 
/* out0172_had-eta12-phi8*/	5, 10, 1, 7, 10, 4, 1, 10, 6, 1, 10, 7, 13, 14, 9, 5, 
/* out0173_had-eta13-phi8*/	4, 14, 8, 6, 14, 9, 11, 14, 10, 7, 14, 11, 1, 
/* out0174_had-eta14-phi8*/	4, 14, 5, 2, 14, 6, 6, 14, 10, 8, 14, 11, 4, 
/* out0175_had-eta15-phi8*/	4, 2, 0, 1, 14, 4, 6, 14, 5, 8, 14, 6, 1, 
/* out0176_had-eta16-phi8*/	2, 2, 0, 12, 14, 4, 1, 
/* out0177_had-eta17-phi8*/	2, 2, 0, 2, 2, 1, 9, 
/* out0178_had-eta18-phi8*/	2, 2, 1, 5, 2, 7, 4, 
/* out0179_had-eta19-phi8*/	1, 2, 7, 1, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 133, 0, 4, 
/* out0182_had-eta2-phi9*/	1, 133, 0, 4, 
/* out0183_had-eta3-phi9*/	5, 104, 0, 8, 105, 2, 4, 106, 0, 7, 106, 1, 15, 132, 0, 5, 
/* out0184_had-eta4-phi9*/	8, 103, 0, 3, 103, 2, 6, 104, 0, 8, 104, 1, 8, 105, 1, 2, 105, 2, 5, 131, 0, 1, 132, 0, 3, 
/* out0185_had-eta5-phi9*/	5, 102, 0, 2, 103, 0, 3, 103, 1, 11, 103, 2, 10, 131, 0, 4, 
/* out0186_had-eta6-phi9*/	6, 64, 2, 3, 102, 0, 14, 102, 1, 4, 103, 1, 1, 130, 0, 1, 131, 0, 3, 
/* out0187_had-eta7-phi9*/	4, 63, 0, 2, 63, 2, 12, 102, 1, 5, 130, 0, 3, 
/* out0188_had-eta8-phi9*/	4, 62, 0, 2, 63, 1, 8, 63, 2, 4, 130, 0, 3, 
/* out0189_had-eta9-phi9*/	4, 62, 0, 11, 62, 1, 1, 129, 0, 3, 130, 0, 1, 
/* out0190_had-eta10-phi9*/	5, 15, 8, 3, 15, 9, 6, 62, 0, 1, 62, 1, 7, 129, 0, 5, 
/* out0191_had-eta11-phi9*/	4, 15, 8, 13, 15, 9, 4, 15, 10, 8, 15, 11, 9, 
/* out0192_had-eta12-phi9*/	5, 14, 3, 5, 15, 4, 1, 15, 5, 13, 15, 6, 1, 15, 11, 7, 
/* out0193_had-eta13-phi9*/	5, 14, 0, 4, 14, 1, 1, 14, 2, 8, 14, 3, 11, 14, 10, 1, 
/* out0194_had-eta14-phi9*/	4, 14, 1, 2, 14, 2, 8, 14, 6, 8, 14, 7, 2, 
/* out0195_had-eta15-phi9*/	4, 14, 4, 8, 14, 6, 1, 14, 7, 7, 18, 8, 1, 
/* out0196_had-eta16-phi9*/	2, 14, 4, 1, 18, 8, 12, 
/* out0197_had-eta17-phi9*/	2, 18, 8, 2, 18, 11, 9, 
/* out0198_had-eta18-phi9*/	2, 18, 5, 4, 18, 11, 5, 
/* out0199_had-eta19-phi9*/	1, 18, 5, 1, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 133, 0, 4, 
/* out0202_had-eta2-phi10*/	4, 106, 0, 2, 107, 0, 4, 107, 2, 8, 133, 0, 4, 
/* out0203_had-eta3-phi10*/	9, 66, 2, 1, 105, 0, 10, 105, 2, 5, 106, 0, 7, 106, 1, 1, 107, 0, 1, 107, 1, 11, 107, 2, 8, 132, 0, 5, 
/* out0204_had-eta4-phi10*/	7, 65, 2, 6, 103, 0, 3, 105, 0, 6, 105, 1, 14, 105, 2, 2, 131, 0, 1, 132, 0, 3, 
/* out0205_had-eta5-phi10*/	7, 64, 0, 3, 64, 2, 3, 65, 1, 3, 65, 2, 7, 103, 0, 7, 103, 1, 4, 131, 0, 4, 
/* out0206_had-eta6-phi10*/	5, 64, 0, 5, 64, 1, 7, 64, 2, 10, 130, 0, 1, 131, 0, 3, 
/* out0207_had-eta7-phi10*/	4, 63, 0, 11, 64, 1, 5, 75, 2, 2, 130, 0, 3, 
/* out0208_had-eta8-phi10*/	4, 63, 0, 3, 63, 1, 8, 74, 2, 3, 130, 0, 3, 
/* out0209_had-eta9-phi10*/	5, 62, 0, 1, 74, 1, 1, 74, 2, 11, 129, 0, 3, 130, 0, 1, 
/* out0210_had-eta10-phi10*/	7, 15, 0, 2, 15, 3, 13, 15, 9, 5, 62, 0, 1, 74, 1, 3, 74, 2, 1, 129, 0, 5, 
/* out0211_had-eta11-phi10*/	7, 15, 0, 1, 15, 1, 1, 15, 2, 16, 15, 3, 3, 15, 6, 6, 15, 9, 1, 15, 10, 8, 
/* out0212_had-eta12-phi10*/	4, 15, 4, 11, 15, 5, 3, 15, 6, 9, 15, 7, 6, 
/* out0213_had-eta13-phi10*/	3, 14, 0, 11, 15, 4, 3, 19, 8, 9, 
/* out0214_had-eta14-phi10*/	4, 14, 0, 1, 14, 1, 13, 14, 7, 1, 19, 11, 5, 
/* out0215_had-eta15-phi10*/	3, 14, 7, 6, 18, 3, 2, 18, 9, 9, 
/* out0216_had-eta16-phi10*/	3, 18, 8, 1, 18, 9, 7, 18, 10, 6, 
/* out0217_had-eta17-phi10*/	3, 18, 6, 2, 18, 10, 8, 18, 11, 2, 
/* out0218_had-eta18-phi10*/	2, 18, 5, 8, 18, 6, 2, 
/* out0219_had-eta19-phi10*/	2, 18, 4, 2, 18, 5, 2, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 138, 0, 4, 
/* out0222_had-eta2-phi11*/	4, 67, 0, 1, 67, 1, 12, 107, 0, 7, 138, 0, 4, 
/* out0223_had-eta3-phi11*/	8, 66, 0, 11, 66, 1, 1, 66, 2, 12, 67, 0, 6, 67, 1, 4, 107, 0, 4, 107, 1, 5, 137, 0, 5, 
/* out0224_had-eta4-phi11*/	7, 65, 0, 11, 65, 2, 2, 66, 1, 13, 66, 2, 3, 77, 2, 3, 136, 0, 1, 137, 0, 3, 
/* out0225_had-eta5-phi11*/	6, 64, 0, 1, 65, 0, 5, 65, 1, 13, 65, 2, 1, 76, 2, 6, 136, 0, 4, 
/* out0226_had-eta6-phi11*/	8, 64, 0, 7, 64, 1, 3, 75, 0, 1, 75, 2, 1, 76, 1, 3, 76, 2, 8, 135, 0, 1, 136, 0, 3, 
/* out0227_had-eta7-phi11*/	5, 64, 1, 1, 75, 0, 4, 75, 1, 2, 75, 2, 11, 135, 0, 3, 
/* out0228_had-eta8-phi11*/	4, 74, 0, 6, 75, 1, 7, 75, 2, 2, 135, 0, 3, 
/* out0229_had-eta9-phi11*/	5, 74, 0, 7, 74, 1, 4, 74, 2, 1, 134, 0, 3, 135, 0, 1, 
/* out0230_had-eta10-phi11*/	4, 15, 0, 5, 20, 2, 3, 74, 1, 7, 134, 0, 5, 
/* out0231_had-eta11-phi11*/	3, 15, 0, 8, 15, 1, 13, 20, 2, 3, 
/* out0232_had-eta12-phi11*/	6, 15, 1, 2, 15, 4, 1, 15, 7, 10, 19, 3, 2, 19, 8, 1, 19, 9, 11, 
/* out0233_had-eta13-phi11*/	4, 19, 8, 6, 19, 9, 5, 19, 10, 10, 19, 11, 3, 
/* out0234_had-eta14-phi11*/	4, 19, 5, 7, 19, 6, 3, 19, 10, 3, 19, 11, 8, 
/* out0235_had-eta15-phi11*/	3, 18, 0, 1, 18, 3, 10, 19, 5, 5, 
/* out0236_had-eta16-phi11*/	3, 18, 2, 9, 18, 3, 4, 18, 10, 1, 
/* out0237_had-eta17-phi11*/	3, 18, 2, 4, 18, 6, 7, 18, 10, 1, 
/* out0238_had-eta18-phi11*/	4, 18, 4, 3, 18, 5, 1, 18, 6, 4, 18, 7, 2, 
/* out0239_had-eta19-phi11*/	1, 18, 4, 7, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 138, 0, 4, 
/* out0242_had-eta2-phi12*/	2, 67, 0, 2, 138, 0, 4, 
/* out0243_had-eta3-phi12*/	6, 66, 0, 4, 67, 0, 7, 78, 0, 7, 78, 1, 6, 78, 2, 16, 137, 0, 5, 
/* out0244_had-eta4-phi12*/	8, 66, 0, 1, 66, 1, 2, 77, 0, 12, 77, 1, 3, 77, 2, 11, 78, 1, 4, 136, 0, 1, 137, 0, 3, 
/* out0245_had-eta5-phi12*/	6, 76, 0, 11, 76, 2, 1, 77, 1, 11, 77, 2, 2, 86, 2, 2, 136, 0, 4, 
/* out0246_had-eta6-phi12*/	7, 75, 0, 1, 76, 0, 4, 76, 1, 13, 76, 2, 1, 85, 2, 3, 135, 0, 1, 136, 0, 3, 
/* out0247_had-eta7-phi12*/	4, 75, 0, 10, 75, 1, 2, 85, 2, 6, 135, 0, 3, 
/* out0248_had-eta8-phi12*/	4, 75, 1, 5, 84, 0, 1, 84, 2, 9, 135, 0, 3, 
/* out0249_had-eta9-phi12*/	6, 74, 0, 3, 74, 1, 1, 84, 1, 3, 84, 2, 6, 134, 0, 3, 135, 0, 1, 
/* out0250_had-eta10-phi12*/	3, 20, 0, 4, 20, 2, 6, 134, 0, 5, 
/* out0251_had-eta11-phi12*/	2, 20, 1, 4, 20, 2, 4, 
/* out0252_had-eta12-phi12*/	3, 19, 0, 5, 19, 3, 12, 20, 1, 3, 
/* out0253_had-eta13-phi12*/	6, 19, 0, 1, 19, 1, 1, 19, 2, 16, 19, 3, 2, 19, 6, 2, 19, 10, 3, 
/* out0254_had-eta14-phi12*/	4, 19, 4, 3, 19, 5, 3, 19, 6, 11, 19, 7, 3, 
/* out0255_had-eta15-phi12*/	4, 6, 8, 1, 18, 0, 6, 19, 4, 10, 19, 5, 1, 
/* out0256_had-eta16-phi12*/	3, 18, 0, 8, 18, 1, 5, 18, 2, 1, 
/* out0257_had-eta17-phi12*/	4, 18, 1, 6, 18, 2, 2, 18, 6, 1, 18, 7, 3, 
/* out0258_had-eta18-phi12*/	2, 18, 4, 2, 18, 7, 8, 
/* out0259_had-eta19-phi12*/	2, 4, 4, 14, 18, 4, 2, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 143, 0, 4, 
/* out0262_had-eta2-phi13*/	1, 143, 0, 4, 
/* out0263_had-eta3-phi13*/	7, 78, 0, 9, 78, 1, 5, 87, 0, 4, 87, 2, 2, 88, 0, 6, 88, 1, 16, 142, 0, 5, 
/* out0264_had-eta4-phi13*/	9, 77, 0, 4, 77, 1, 1, 78, 1, 1, 86, 0, 1, 87, 0, 3, 87, 1, 8, 87, 2, 14, 141, 0, 1, 142, 0, 3, 
/* out0265_had-eta5-phi13*/	5, 77, 1, 1, 86, 0, 8, 86, 1, 4, 86, 2, 13, 141, 0, 4, 
/* out0266_had-eta6-phi13*/	7, 76, 0, 1, 85, 0, 10, 85, 2, 3, 86, 1, 7, 86, 2, 1, 140, 0, 1, 141, 0, 3, 
/* out0267_had-eta7-phi13*/	4, 85, 0, 2, 85, 1, 12, 85, 2, 4, 140, 0, 3, 
/* out0268_had-eta8-phi13*/	4, 84, 0, 13, 84, 2, 1, 85, 1, 1, 140, 0, 3, 
/* out0269_had-eta9-phi13*/	3, 84, 1, 11, 139, 0, 3, 140, 0, 1, 
/* out0270_had-eta10-phi13*/	3, 20, 0, 9, 28, 2, 1, 139, 0, 5, 
/* out0271_had-eta11-phi13*/	3, 7, 9, 1, 20, 0, 2, 20, 1, 6, 
/* out0272_had-eta12-phi13*/	3, 7, 8, 12, 19, 0, 6, 20, 1, 2, 
/* out0273_had-eta13-phi13*/	4, 7, 8, 2, 7, 11, 4, 19, 0, 4, 19, 1, 14, 
/* out0274_had-eta14-phi13*/	4, 6, 9, 4, 19, 1, 1, 19, 4, 1, 19, 7, 13, 
/* out0275_had-eta15-phi13*/	3, 6, 8, 11, 6, 9, 4, 19, 4, 2, 
/* out0276_had-eta16-phi13*/	4, 6, 8, 4, 6, 11, 7, 18, 0, 1, 18, 1, 1, 
/* out0277_had-eta17-phi13*/	4, 6, 5, 1, 6, 11, 4, 18, 1, 4, 18, 7, 1, 
/* out0278_had-eta18-phi13*/	2, 4, 5, 8, 18, 7, 2, 
/* out0279_had-eta19-phi13*/	3, 4, 4, 2, 4, 5, 6, 4, 6, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 143, 0, 4, 
/* out0282_had-eta2-phi14*/	1, 143, 0, 4, 
/* out0283_had-eta3-phi14*/	3, 87, 0, 3, 88, 0, 10, 142, 0, 5, 
/* out0284_had-eta4-phi14*/	6, 31, 0, 4, 31, 2, 8, 87, 0, 6, 87, 1, 8, 141, 0, 1, 142, 0, 3, 
/* out0285_had-eta5-phi14*/	7, 30, 0, 2, 30, 2, 1, 31, 1, 4, 31, 2, 8, 86, 0, 7, 86, 1, 3, 141, 0, 4, 
/* out0286_had-eta6-phi14*/	7, 30, 0, 1, 30, 1, 2, 30, 2, 14, 85, 0, 2, 86, 1, 2, 140, 0, 1, 141, 0, 3, 
/* out0287_had-eta7-phi14*/	7, 29, 0, 4, 29, 2, 6, 30, 1, 2, 30, 2, 1, 85, 0, 2, 85, 1, 3, 140, 0, 3, 
/* out0288_had-eta8-phi14*/	4, 29, 1, 3, 29, 2, 10, 84, 0, 2, 140, 0, 3, 
/* out0289_had-eta9-phi14*/	6, 28, 0, 4, 28, 2, 6, 29, 1, 1, 84, 1, 2, 139, 0, 3, 140, 0, 1, 
/* out0290_had-eta10-phi14*/	3, 28, 1, 2, 28, 2, 8, 139, 0, 5, 
/* out0291_had-eta11-phi14*/	6, 7, 3, 12, 7, 9, 8, 20, 0, 1, 20, 1, 1, 28, 1, 2, 28, 2, 1, 
/* out0292_had-eta12-phi14*/	6, 7, 2, 3, 7, 6, 1, 7, 8, 2, 7, 9, 7, 7, 10, 14, 7, 11, 2, 
/* out0293_had-eta13-phi14*/	4, 7, 5, 9, 7, 6, 3, 7, 10, 2, 7, 11, 10, 
/* out0294_had-eta14-phi14*/	3, 6, 3, 12, 6, 9, 5, 7, 5, 3, 
/* out0295_had-eta15-phi14*/	3, 6, 2, 4, 6, 9, 3, 6, 10, 10, 
/* out0296_had-eta16-phi14*/	4, 6, 5, 1, 6, 6, 4, 6, 10, 6, 6, 11, 4, 
/* out0297_had-eta17-phi14*/	3, 4, 3, 1, 6, 5, 10, 6, 11, 1, 
/* out0298_had-eta18-phi14*/	2, 4, 3, 9, 4, 5, 1, 
/* out0299_had-eta19-phi14*/	4, 4, 2, 5, 4, 3, 1, 4, 5, 1, 4, 6, 15, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 148, 0, 4, 
/* out0302_had-eta2-phi15*/	1, 148, 0, 4, 
/* out0303_had-eta3-phi15*/	5, 40, 0, 2, 40, 2, 1, 41, 0, 2, 41, 1, 16, 147, 0, 5, 
/* out0304_had-eta4-phi15*/	5, 31, 0, 12, 40, 1, 1, 40, 2, 13, 146, 0, 1, 147, 0, 3, 
/* out0305_had-eta5-phi15*/	5, 30, 0, 4, 31, 1, 12, 39, 0, 1, 39, 2, 9, 146, 0, 4, 
/* out0306_had-eta6-phi15*/	6, 30, 0, 9, 30, 1, 9, 38, 2, 2, 39, 2, 2, 145, 0, 1, 146, 0, 3, 
/* out0307_had-eta7-phi15*/	4, 29, 0, 10, 30, 1, 3, 38, 2, 5, 145, 0, 3, 
/* out0308_had-eta8-phi15*/	4, 29, 0, 2, 29, 1, 11, 37, 2, 1, 145, 0, 3, 
/* out0309_had-eta9-phi15*/	5, 28, 0, 10, 29, 1, 1, 37, 2, 2, 144, 0, 3, 145, 0, 1, 
/* out0310_had-eta10-phi15*/	3, 28, 0, 2, 28, 1, 9, 144, 0, 5, 
/* out0311_had-eta11-phi15*/	6, 7, 0, 15, 7, 1, 1, 7, 2, 1, 7, 3, 4, 13, 2, 1, 28, 1, 2, 
/* out0312_had-eta12-phi15*/	4, 7, 1, 7, 7, 2, 12, 7, 6, 7, 7, 7, 3, 
/* out0313_had-eta13-phi15*/	4, 7, 4, 11, 7, 5, 4, 7, 6, 5, 7, 7, 4, 
/* out0314_had-eta14-phi15*/	3, 6, 0, 12, 6, 3, 4, 7, 4, 2, 
/* out0315_had-eta15-phi15*/	3, 6, 1, 3, 6, 2, 12, 6, 6, 2, 
/* out0316_had-eta16-phi15*/	4, 6, 4, 1, 6, 5, 1, 6, 6, 10, 6, 7, 2, 
/* out0317_had-eta17-phi15*/	3, 4, 0, 1, 6, 4, 8, 6, 5, 3, 
/* out0318_had-eta18-phi15*/	2, 4, 0, 6, 4, 3, 4, 
/* out0319_had-eta19-phi15*/	3, 4, 1, 1, 4, 2, 10, 4, 3, 1, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 148, 0, 4, 
/* out0322_had-eta2-phi16*/	1, 148, 0, 4, 
/* out0323_had-eta3-phi16*/	5, 40, 0, 6, 41, 0, 14, 51, 0, 2, 51, 2, 13, 147, 0, 5, 
/* out0324_had-eta4-phi16*/	8, 39, 0, 1, 40, 0, 8, 40, 1, 15, 40, 2, 2, 50, 2, 5, 51, 2, 1, 146, 0, 1, 147, 0, 3, 
/* out0325_had-eta5-phi16*/	5, 39, 0, 14, 39, 1, 7, 39, 2, 4, 50, 2, 1, 146, 0, 4, 
/* out0326_had-eta6-phi16*/	7, 38, 0, 11, 38, 2, 2, 39, 1, 8, 39, 2, 1, 49, 2, 1, 145, 0, 1, 146, 0, 3, 
/* out0327_had-eta7-phi16*/	4, 38, 0, 2, 38, 1, 10, 38, 2, 7, 145, 0, 3, 
/* out0328_had-eta8-phi16*/	4, 37, 0, 8, 37, 2, 6, 38, 1, 1, 145, 0, 3, 
/* out0329_had-eta9-phi16*/	4, 37, 1, 5, 37, 2, 7, 144, 0, 3, 145, 0, 1, 
/* out0330_had-eta10-phi16*/	4, 13, 0, 3, 13, 2, 5, 28, 1, 1, 144, 0, 5, 
/* out0331_had-eta11-phi16*/	2, 7, 0, 1, 13, 2, 8, 
/* out0332_had-eta12-phi16*/	6, 7, 1, 8, 7, 7, 6, 11, 3, 2, 11, 9, 4, 13, 1, 1, 13, 2, 1, 
/* out0333_had-eta13-phi16*/	5, 7, 4, 3, 7, 7, 3, 11, 8, 7, 11, 9, 11, 11, 10, 1, 
/* out0334_had-eta14-phi16*/	4, 6, 0, 4, 6, 1, 1, 11, 8, 9, 11, 11, 6, 
/* out0335_had-eta15-phi16*/	3, 6, 1, 12, 6, 7, 3, 11, 11, 2, 
/* out0336_had-eta16-phi16*/	4, 5, 8, 1, 5, 9, 1, 6, 4, 2, 6, 7, 10, 
/* out0337_had-eta17-phi16*/	3, 4, 0, 1, 5, 8, 6, 6, 4, 5, 
/* out0338_had-eta18-phi16*/	2, 4, 0, 8, 5, 8, 2, 
/* out0339_had-eta19-phi16*/	2, 4, 1, 10, 4, 2, 1, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 153, 0, 4, 
/* out0342_had-eta2-phi17*/	2, 61, 1, 5, 153, 0, 4, 
/* out0343_had-eta3-phi17*/	7, 51, 0, 14, 51, 1, 12, 51, 2, 2, 60, 2, 4, 61, 0, 1, 61, 1, 11, 152, 0, 5, 
/* out0344_had-eta4-phi17*/	7, 50, 0, 15, 50, 1, 5, 50, 2, 6, 51, 1, 4, 60, 2, 3, 151, 0, 1, 152, 0, 3, 
/* out0345_had-eta5-phi17*/	6, 39, 1, 1, 49, 0, 9, 49, 2, 3, 50, 1, 9, 50, 2, 4, 151, 0, 4, 
/* out0346_had-eta6-phi17*/	6, 38, 0, 2, 49, 0, 1, 49, 1, 6, 49, 2, 12, 150, 0, 1, 151, 0, 3, 
/* out0347_had-eta7-phi17*/	5, 38, 0, 1, 38, 1, 5, 48, 0, 3, 48, 2, 9, 150, 0, 3, 
/* out0348_had-eta8-phi17*/	4, 37, 0, 8, 37, 1, 2, 48, 2, 5, 150, 0, 3, 
/* out0349_had-eta9-phi17*/	5, 13, 0, 1, 37, 1, 9, 47, 2, 3, 149, 0, 3, 150, 0, 1, 
/* out0350_had-eta10-phi17*/	3, 13, 0, 10, 47, 2, 1, 149, 0, 5, 
/* out0351_had-eta11-phi17*/	2, 13, 1, 8, 13, 2, 1, 
/* out0352_had-eta12-phi17*/	3, 11, 0, 6, 11, 3, 12, 13, 1, 3, 
/* out0353_had-eta13-phi17*/	5, 11, 2, 10, 11, 3, 2, 11, 6, 1, 11, 9, 1, 11, 10, 9, 
/* out0354_had-eta14-phi17*/	4, 11, 5, 4, 11, 6, 5, 11, 10, 6, 11, 11, 5, 
/* out0355_had-eta15-phi17*/	5, 5, 3, 5, 5, 9, 1, 6, 7, 1, 11, 5, 7, 11, 11, 3, 
/* out0356_had-eta16-phi17*/	3, 5, 3, 2, 5, 9, 11, 5, 10, 1, 
/* out0357_had-eta17-phi17*/	4, 5, 8, 4, 5, 9, 3, 5, 10, 3, 5, 11, 1, 
/* out0358_had-eta18-phi17*/	2, 5, 8, 3, 5, 11, 7, 
/* out0359_had-eta19-phi17*/	2, 4, 1, 5, 5, 11, 2, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 153, 0, 4, 
/* out0362_had-eta2-phi18*/	4, 61, 0, 7, 101, 0, 3, 101, 2, 4, 153, 0, 4, 
/* out0363_had-eta3-phi18*/	6, 60, 0, 16, 60, 1, 4, 60, 2, 4, 61, 0, 8, 101, 2, 8, 152, 0, 5, 
/* out0364_had-eta4-phi18*/	8, 50, 0, 1, 50, 1, 2, 59, 0, 10, 59, 2, 3, 60, 1, 11, 60, 2, 5, 151, 0, 1, 152, 0, 3, 
/* out0365_had-eta5-phi18*/	6, 49, 0, 6, 58, 0, 1, 59, 0, 1, 59, 1, 5, 59, 2, 13, 151, 0, 4, 
/* out0366_had-eta6-phi18*/	6, 48, 0, 2, 49, 1, 10, 58, 0, 1, 58, 2, 9, 150, 0, 1, 151, 0, 3, 
/* out0367_had-eta7-phi18*/	5, 48, 0, 11, 48, 1, 6, 48, 2, 1, 58, 2, 1, 150, 0, 3, 
/* out0368_had-eta8-phi18*/	4, 47, 0, 6, 48, 1, 9, 48, 2, 1, 150, 0, 3, 
/* out0369_had-eta9-phi18*/	5, 47, 0, 3, 47, 1, 1, 47, 2, 8, 149, 0, 3, 150, 0, 1, 
/* out0370_had-eta10-phi18*/	7, 12, 3, 4, 12, 9, 1, 13, 0, 2, 13, 1, 1, 47, 1, 3, 47, 2, 4, 149, 0, 5, 
/* out0371_had-eta11-phi18*/	4, 12, 3, 1, 12, 8, 6, 12, 9, 14, 13, 1, 3, 
/* out0372_had-eta12-phi18*/	4, 11, 0, 10, 11, 1, 4, 12, 8, 10, 12, 11, 3, 
/* out0373_had-eta13-phi18*/	4, 11, 1, 9, 11, 2, 6, 11, 6, 5, 11, 7, 5, 
/* out0374_had-eta14-phi18*/	4, 11, 4, 8, 11, 5, 3, 11, 6, 5, 11, 7, 4, 
/* out0375_had-eta15-phi18*/	4, 5, 0, 6, 5, 3, 5, 11, 4, 4, 11, 5, 2, 
/* out0376_had-eta16-phi18*/	3, 5, 2, 8, 5, 3, 4, 5, 10, 2, 
/* out0377_had-eta17-phi18*/	3, 5, 2, 1, 5, 6, 2, 5, 10, 8, 
/* out0378_had-eta18-phi18*/	4, 5, 5, 3, 5, 6, 2, 5, 10, 2, 5, 11, 4, 
/* out0379_had-eta19-phi18*/	2, 5, 5, 5, 5, 11, 2, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 158, 0, 4, 
/* out0382_had-eta2-phi19*/	4, 100, 1, 1, 101, 0, 13, 101, 1, 2, 158, 0, 4, 
/* out0383_had-eta3-phi19*/	7, 60, 1, 1, 99, 0, 13, 99, 2, 3, 100, 1, 5, 101, 1, 14, 101, 2, 4, 157, 0, 5, 
/* out0384_had-eta4-phi19*/	9, 59, 0, 5, 59, 1, 1, 98, 0, 3, 98, 2, 1, 99, 0, 1, 99, 1, 9, 99, 2, 13, 156, 0, 1, 157, 0, 3, 
/* out0385_had-eta5-phi19*/	4, 58, 0, 6, 59, 1, 10, 98, 2, 10, 156, 0, 4, 
/* out0386_had-eta6-phi19*/	5, 58, 0, 8, 58, 1, 10, 58, 2, 4, 155, 0, 1, 156, 0, 3, 
/* out0387_had-eta7-phi19*/	6, 48, 1, 1, 57, 0, 7, 57, 2, 5, 58, 1, 3, 58, 2, 2, 155, 0, 3, 
/* out0388_had-eta8-phi19*/	3, 47, 0, 3, 57, 2, 11, 155, 0, 3, 
/* out0389_had-eta9-phi19*/	5, 47, 0, 4, 47, 1, 8, 68, 2, 1, 154, 0, 3, 155, 0, 1, 
/* out0390_had-eta10-phi19*/	5, 12, 0, 13, 12, 1, 1, 12, 3, 8, 47, 1, 4, 154, 0, 5, 
/* out0391_had-eta11-phi19*/	6, 12, 1, 1, 12, 2, 14, 12, 3, 3, 12, 6, 4, 12, 9, 1, 12, 10, 11, 
/* out0392_had-eta12-phi19*/	4, 12, 5, 8, 12, 6, 4, 12, 10, 5, 12, 11, 12, 
/* out0393_had-eta13-phi19*/	6, 11, 1, 3, 11, 7, 6, 12, 5, 2, 12, 11, 1, 16, 3, 3, 16, 9, 7, 
/* out0394_had-eta14-phi19*/	4, 11, 4, 4, 11, 7, 1, 16, 8, 8, 16, 9, 4, 
/* out0395_had-eta15-phi19*/	3, 5, 0, 9, 5, 1, 1, 16, 8, 5, 
/* out0396_had-eta16-phi19*/	4, 5, 0, 1, 5, 1, 7, 5, 2, 6, 5, 6, 1, 
/* out0397_had-eta17-phi19*/	3, 5, 2, 1, 5, 6, 9, 5, 7, 2, 
/* out0398_had-eta18-phi19*/	3, 5, 4, 2, 5, 5, 5, 5, 6, 2, 
/* out0399_had-eta19-phi19*/	2, 5, 4, 1, 5, 5, 3, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 158, 0, 4, 
/* out0402_had-eta2-phi20*/	1, 158, 0, 4, 
/* out0403_had-eta3-phi20*/	7, 99, 0, 2, 99, 1, 1, 100, 0, 16, 100, 1, 10, 112, 0, 7, 112, 2, 1, 157, 0, 5, 
/* out0404_had-eta4-phi20*/	6, 98, 0, 9, 99, 1, 6, 112, 0, 1, 112, 2, 15, 156, 0, 1, 157, 0, 3, 
/* out0405_had-eta5-phi20*/	5, 98, 0, 4, 98, 1, 16, 98, 2, 5, 108, 0, 2, 156, 0, 4, 
/* out0406_had-eta6-phi20*/	5, 58, 1, 3, 108, 0, 6, 108, 2, 11, 155, 0, 1, 156, 0, 3, 
/* out0407_had-eta7-phi20*/	4, 57, 0, 9, 57, 1, 4, 108, 2, 5, 155, 0, 3, 
/* out0408_had-eta8-phi20*/	3, 57, 1, 12, 68, 0, 2, 155, 0, 3, 
/* out0409_had-eta9-phi20*/	4, 68, 0, 5, 68, 2, 7, 154, 0, 3, 155, 0, 1, 
/* out0410_had-eta10-phi20*/	4, 12, 0, 3, 12, 1, 6, 68, 2, 8, 154, 0, 5, 
/* out0411_had-eta11-phi20*/	5, 12, 1, 8, 12, 2, 2, 12, 4, 2, 12, 6, 6, 12, 7, 16, 
/* out0412_had-eta12-phi20*/	4, 12, 4, 14, 12, 5, 6, 12, 6, 2, 16, 0, 5, 
/* out0413_had-eta13-phi20*/	5, 16, 0, 3, 16, 2, 6, 16, 3, 13, 16, 9, 2, 16, 10, 1, 
/* out0414_had-eta14-phi20*/	5, 16, 2, 1, 16, 8, 1, 16, 9, 3, 16, 10, 13, 16, 11, 1, 
/* out0415_had-eta15-phi20*/	4, 5, 1, 1, 16, 8, 2, 16, 10, 1, 16, 11, 13, 
/* out0416_had-eta16-phi20*/	3, 5, 1, 7, 5, 7, 6, 16, 11, 1, 
/* out0417_had-eta17-phi20*/	2, 5, 4, 3, 5, 7, 8, 
/* out0418_had-eta18-phi20*/	1, 5, 4, 9, 
/* out0419_had-eta19-phi20*/	1, 5, 4, 1, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 163, 0, 4, 
/* out0422_had-eta2-phi21*/	1, 163, 0, 4, 
/* out0423_had-eta3-phi21*/	7, 110, 0, 2, 110, 2, 1, 112, 0, 7, 112, 1, 1, 113, 0, 10, 113, 1, 16, 162, 0, 5, 
/* out0424_had-eta4-phi21*/	6, 109, 0, 9, 110, 2, 6, 112, 0, 1, 112, 1, 15, 161, 0, 1, 162, 0, 3, 
/* out0425_had-eta5-phi21*/	5, 108, 0, 2, 109, 0, 4, 109, 1, 5, 109, 2, 16, 161, 0, 4, 
/* out0426_had-eta6-phi21*/	5, 70, 2, 3, 108, 0, 6, 108, 1, 11, 160, 0, 1, 161, 0, 3, 
/* out0427_had-eta7-phi21*/	4, 69, 0, 9, 69, 2, 4, 108, 1, 5, 160, 0, 3, 
/* out0428_had-eta8-phi21*/	3, 68, 0, 3, 69, 2, 12, 160, 0, 3, 
/* out0429_had-eta9-phi21*/	4, 68, 0, 6, 68, 1, 6, 159, 0, 3, 160, 0, 1, 
/* out0430_had-eta10-phi21*/	4, 17, 0, 3, 17, 3, 6, 68, 1, 8, 159, 0, 5, 
/* out0431_had-eta11-phi21*/	5, 17, 2, 2, 17, 3, 8, 17, 8, 2, 17, 9, 16, 17, 10, 6, 
/* out0432_had-eta12-phi21*/	4, 16, 0, 5, 17, 8, 14, 17, 10, 2, 17, 11, 6, 
/* out0433_had-eta13-phi21*/	5, 16, 0, 3, 16, 1, 12, 16, 2, 7, 16, 6, 1, 16, 7, 1, 
/* out0434_had-eta14-phi21*/	5, 16, 2, 2, 16, 5, 1, 16, 6, 14, 16, 7, 2, 16, 10, 1, 
/* out0435_had-eta15-phi21*/	5, 16, 4, 1, 16, 5, 14, 16, 6, 1, 16, 11, 1, 21, 3, 1, 
/* out0436_had-eta16-phi21*/	3, 16, 5, 1, 21, 3, 7, 21, 9, 6, 
/* out0437_had-eta17-phi21*/	2, 21, 8, 3, 21, 9, 8, 
/* out0438_had-eta18-phi21*/	1, 21, 8, 9, 
/* out0439_had-eta19-phi21*/	1, 21, 8, 1, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 163, 0, 4, 
/* out0442_had-eta2-phi22*/	4, 111, 0, 13, 111, 2, 2, 113, 0, 1, 163, 0, 4, 
/* out0443_had-eta3-phi22*/	7, 72, 2, 1, 110, 0, 13, 110, 1, 3, 111, 1, 4, 111, 2, 14, 113, 0, 5, 162, 0, 5, 
/* out0444_had-eta4-phi22*/	9, 71, 0, 5, 71, 2, 1, 109, 0, 3, 109, 1, 1, 110, 0, 1, 110, 1, 13, 110, 2, 9, 161, 0, 1, 162, 0, 3, 
/* out0445_had-eta5-phi22*/	4, 70, 0, 6, 71, 2, 10, 109, 1, 10, 161, 0, 4, 
/* out0446_had-eta6-phi22*/	5, 70, 0, 8, 70, 1, 4, 70, 2, 10, 160, 0, 1, 161, 0, 3, 
/* out0447_had-eta7-phi22*/	6, 69, 0, 7, 69, 1, 5, 70, 1, 2, 70, 2, 3, 80, 2, 1, 160, 0, 3, 
/* out0448_had-eta8-phi22*/	3, 69, 1, 11, 79, 0, 3, 160, 0, 3, 
/* out0449_had-eta9-phi22*/	5, 68, 1, 1, 79, 0, 4, 79, 2, 8, 159, 0, 3, 160, 0, 1, 
/* out0450_had-eta10-phi22*/	6, 17, 0, 13, 17, 1, 8, 17, 3, 1, 68, 1, 1, 79, 2, 4, 159, 0, 5, 
/* out0451_had-eta11-phi22*/	6, 17, 1, 3, 17, 2, 14, 17, 3, 1, 17, 6, 11, 17, 7, 1, 17, 10, 4, 
/* out0452_had-eta12-phi22*/	4, 17, 5, 12, 17, 6, 5, 17, 10, 4, 17, 11, 8, 
/* out0453_had-eta13-phi22*/	6, 16, 1, 4, 16, 7, 8, 17, 5, 1, 17, 11, 2, 22, 3, 3, 22, 9, 6, 
/* out0454_had-eta14-phi22*/	4, 16, 4, 9, 16, 7, 5, 22, 8, 4, 22, 9, 1, 
/* out0455_had-eta15-phi22*/	3, 16, 4, 6, 21, 0, 9, 21, 3, 1, 
/* out0456_had-eta16-phi22*/	4, 21, 0, 1, 21, 2, 6, 21, 3, 7, 21, 10, 1, 
/* out0457_had-eta17-phi22*/	3, 21, 2, 1, 21, 9, 2, 21, 10, 9, 
/* out0458_had-eta18-phi22*/	3, 21, 8, 2, 21, 10, 2, 21, 11, 5, 
/* out0459_had-eta19-phi22*/	2, 21, 8, 1, 21, 11, 3, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 168, 0, 4, 
/* out0462_had-eta2-phi23*/	4, 73, 1, 7, 111, 0, 3, 111, 1, 4, 168, 0, 4, 
/* out0463_had-eta3-phi23*/	6, 72, 0, 16, 72, 1, 4, 72, 2, 4, 73, 1, 8, 111, 1, 8, 167, 0, 5, 
/* out0464_had-eta4-phi23*/	8, 71, 0, 10, 71, 1, 3, 72, 1, 5, 72, 2, 11, 82, 0, 1, 82, 2, 2, 166, 0, 1, 167, 0, 3, 
/* out0465_had-eta5-phi23*/	6, 70, 0, 1, 71, 0, 1, 71, 1, 13, 71, 2, 5, 81, 0, 6, 166, 0, 4, 
/* out0466_had-eta6-phi23*/	6, 70, 0, 1, 70, 1, 9, 80, 0, 2, 81, 2, 10, 165, 0, 1, 166, 0, 3, 
/* out0467_had-eta7-phi23*/	5, 70, 1, 1, 80, 0, 11, 80, 1, 1, 80, 2, 6, 165, 0, 3, 
/* out0468_had-eta8-phi23*/	4, 79, 0, 6, 80, 1, 1, 80, 2, 9, 165, 0, 3, 
/* out0469_had-eta9-phi23*/	5, 79, 0, 3, 79, 1, 8, 79, 2, 1, 164, 0, 3, 165, 0, 1, 
/* out0470_had-eta10-phi23*/	7, 17, 1, 4, 17, 7, 1, 23, 0, 2, 23, 2, 1, 79, 1, 4, 79, 2, 3, 164, 0, 5, 
/* out0471_had-eta11-phi23*/	4, 17, 1, 1, 17, 4, 6, 17, 7, 14, 23, 2, 3, 
/* out0472_had-eta12-phi23*/	4, 17, 4, 10, 17, 5, 3, 22, 0, 10, 22, 3, 4, 
/* out0473_had-eta13-phi23*/	4, 22, 2, 6, 22, 3, 9, 22, 9, 5, 22, 10, 5, 
/* out0474_had-eta14-phi23*/	4, 22, 8, 8, 22, 9, 4, 22, 10, 5, 22, 11, 3, 
/* out0475_had-eta15-phi23*/	4, 21, 0, 6, 21, 1, 5, 22, 8, 4, 22, 11, 2, 
/* out0476_had-eta16-phi23*/	3, 21, 1, 4, 21, 2, 8, 21, 6, 2, 
/* out0477_had-eta17-phi23*/	3, 21, 2, 1, 21, 6, 8, 21, 10, 2, 
/* out0478_had-eta18-phi23*/	4, 21, 5, 4, 21, 6, 2, 21, 10, 2, 21, 11, 3, 
/* out0479_had-eta19-phi23*/	2, 21, 5, 2, 21, 11, 5, 
/* out0480_had-eta0-phi24*/	0, 
/* out0481_had-eta1-phi24*/	1, 168, 0, 4, 
/* out0482_had-eta2-phi24*/	2, 73, 0, 5, 168, 0, 4, 
/* out0483_had-eta3-phi24*/	7, 72, 1, 4, 73, 0, 11, 73, 1, 1, 83, 0, 14, 83, 1, 2, 83, 2, 12, 167, 0, 5, 
/* out0484_had-eta4-phi24*/	7, 72, 1, 3, 82, 0, 15, 82, 1, 6, 82, 2, 5, 83, 2, 4, 166, 0, 1, 167, 0, 3, 
/* out0485_had-eta5-phi24*/	6, 81, 0, 9, 81, 1, 3, 82, 1, 4, 82, 2, 9, 91, 2, 1, 166, 0, 4, 
/* out0486_had-eta6-phi24*/	6, 81, 0, 1, 81, 1, 12, 81, 2, 6, 90, 0, 3, 165, 0, 1, 166, 0, 3, 
/* out0487_had-eta7-phi24*/	5, 80, 0, 3, 80, 1, 9, 90, 0, 1, 90, 2, 5, 165, 0, 3, 
/* out0488_had-eta8-phi24*/	4, 80, 1, 5, 89, 0, 8, 89, 2, 2, 165, 0, 3, 
/* out0489_had-eta9-phi24*/	5, 23, 0, 1, 79, 1, 3, 89, 2, 9, 164, 0, 3, 165, 0, 1, 
/* out0490_had-eta10-phi24*/	3, 23, 0, 10, 79, 1, 1, 164, 0, 5, 
/* out0491_had-eta11-phi24*/	2, 23, 1, 1, 23, 2, 8, 
/* out0492_had-eta12-phi24*/	3, 22, 0, 6, 22, 1, 12, 23, 2, 3, 
/* out0493_had-eta13-phi24*/	5, 22, 1, 2, 22, 2, 10, 22, 6, 9, 22, 7, 1, 22, 10, 1, 
/* out0494_had-eta14-phi24*/	4, 22, 5, 5, 22, 6, 6, 22, 10, 5, 22, 11, 4, 
/* out0495_had-eta15-phi24*/	4, 21, 1, 5, 21, 7, 1, 22, 5, 3, 22, 11, 7, 
/* out0496_had-eta16-phi24*/	3, 21, 1, 2, 21, 6, 1, 21, 7, 11, 
/* out0497_had-eta17-phi24*/	4, 21, 4, 4, 21, 5, 1, 21, 6, 3, 21, 7, 3, 
/* out0498_had-eta18-phi24*/	2, 21, 4, 3, 21, 5, 7, 
/* out0499_had-eta19-phi24*/	1, 21, 5, 2, 
/* out0500_had-eta0-phi25*/	0, 
/* out0501_had-eta1-phi25*/	1, 173, 0, 4, 
/* out0502_had-eta2-phi25*/	1, 173, 0, 4, 
/* out0503_had-eta3-phi25*/	5, 83, 0, 2, 83, 1, 13, 92, 0, 6, 93, 1, 14, 172, 0, 5, 
/* out0504_had-eta4-phi25*/	8, 82, 1, 5, 83, 1, 1, 91, 0, 1, 92, 0, 8, 92, 1, 2, 92, 2, 15, 171, 0, 1, 172, 0, 3, 
/* out0505_had-eta5-phi25*/	5, 82, 1, 1, 91, 0, 14, 91, 1, 4, 91, 2, 7, 171, 0, 4, 
/* out0506_had-eta6-phi25*/	7, 81, 1, 1, 90, 0, 11, 90, 1, 2, 91, 1, 1, 91, 2, 8, 170, 0, 1, 171, 0, 3, 
/* out0507_had-eta7-phi25*/	4, 90, 0, 1, 90, 1, 7, 90, 2, 10, 170, 0, 3, 
/* out0508_had-eta8-phi25*/	4, 89, 0, 8, 89, 1, 6, 90, 2, 1, 170, 0, 3, 
/* out0509_had-eta9-phi25*/	4, 89, 1, 7, 89, 2, 5, 169, 0, 3, 170, 0, 1, 
/* out0510_had-eta10-phi25*/	3, 23, 0, 3, 23, 1, 5, 169, 0, 5, 
/* out0511_had-eta11-phi25*/	1, 23, 1, 8, 
/* out0512_had-eta12-phi25*/	4, 22, 1, 2, 22, 7, 4, 23, 1, 1, 23, 2, 1, 
/* out0513_had-eta13-phi25*/	3, 22, 4, 7, 22, 6, 1, 22, 7, 11, 
/* out0514_had-eta14-phi25*/	2, 22, 4, 9, 22, 5, 6, 
/* out0515_had-eta15-phi25*/	1, 22, 5, 2, 
/* out0516_had-eta16-phi25*/	2, 21, 4, 1, 21, 7, 1, 
/* out0517_had-eta17-phi25*/	1, 21, 4, 6, 
/* out0518_had-eta18-phi25*/	1, 21, 4, 2, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	0, 
/* out0521_had-eta1-phi26*/	1, 173, 0, 4, 
/* out0522_had-eta2-phi26*/	1, 173, 0, 4, 
/* out0523_had-eta3-phi26*/	5, 92, 0, 2, 92, 1, 1, 93, 0, 16, 93, 1, 2, 172, 0, 5, 
/* out0524_had-eta4-phi26*/	4, 92, 1, 13, 92, 2, 1, 171, 0, 1, 172, 0, 3, 
/* out0525_had-eta5-phi26*/	3, 91, 0, 1, 91, 1, 9, 171, 0, 4, 
/* out0526_had-eta6-phi26*/	4, 90, 1, 2, 91, 1, 2, 170, 0, 1, 171, 0, 3, 
/* out0527_had-eta7-phi26*/	2, 90, 1, 5, 170, 0, 3, 
/* out0528_had-eta8-phi26*/	2, 89, 1, 1, 170, 0, 3, 
/* out0529_had-eta9-phi26*/	3, 89, 1, 2, 169, 0, 3, 170, 0, 1, 
/* out0530_had-eta10-phi26*/	1, 169, 0, 5, 
/* out0531_had-eta11-phi26*/	1, 23, 1, 1, 
/* out0532_had-eta12-phi26*/	0, 
/* out0533_had-eta13-phi26*/	0, 
/* out0534_had-eta14-phi26*/	0, 
/* out0535_had-eta15-phi26*/	0, 
/* out0536_had-eta16-phi26*/	0, 
/* out0537_had-eta17-phi26*/	0, 
/* out0538_had-eta18-phi26*/	0, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	0, 
/* out0550_had-eta10-phi27*/	0, 
/* out0551_had-eta11-phi27*/	0, 
/* out0552_had-eta12-phi27*/	0, 
/* out0553_had-eta13-phi27*/	0, 
/* out0554_had-eta14-phi27*/	0, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	0, 
/* out0557_had-eta17-phi27*/	0, 
/* out0558_had-eta18-phi27*/	0, 
/* out0559_had-eta19-phi27*/	0, 
};