parameter integer matrixH [0:8753] = {
/* num inputs = 194(in0-in193) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2757 */

/* out0000_em-eta0-phi0*/	1,149,0,6,
/* out0001_em-eta1-phi0*/	2,148,0,3,149,0,10,
/* out0002_em-eta2-phi0*/	2,148,0,13,148,1,5,
/* out0003_em-eta3-phi0*/	4,60,0,14,60,1,4,147,0,6,148,1,11,
/* out0004_em-eta4-phi0*/	7,51,1,5,59,0,10,59,1,2,60,0,2,60,2,2,147,0,10,147,1,7,
/* out0005_em-eta5-phi0*/	9,51,0,16,51,1,11,51,2,9,58,0,3,58,1,1,59,0,5,59,2,1,146,0,8,147,1,9,
/* out0006_em-eta6-phi0*/	8,50,0,15,50,1,13,50,2,3,51,2,7,58,0,8,63,2,1,146,0,8,146,1,16,
/* out0007_em-eta7-phi0*/	9,49,1,2,50,0,1,50,1,3,50,2,13,57,0,6,62,0,1,62,1,4,63,1,6,63,2,12,
/* out0008_em-eta8-phi0*/	7,49,0,16,49,1,11,49,2,5,57,0,1,62,0,14,62,1,2,62,2,2,
/* out0009_em-eta9-phi0*/	7,48,1,4,49,2,8,56,0,3,61,0,6,61,1,3,62,0,1,62,2,2,
/* out0010_em-eta10-phi0*/	5,48,0,16,48,1,11,48,2,6,61,0,10,61,2,2,
/* out0011_em-eta11-phi0*/	7,7,2,16,7,3,3,18,5,1,19,5,2,48,2,8,60,0,5,60,1,2,
/* out0012_em-eta12-phi0*/	6,6,2,4,6,3,13,7,3,13,7,4,4,18,5,1,60,0,8,
/* out0013_em-eta13-phi0*/	11,6,0,1,6,1,7,6,2,12,6,3,1,7,0,16,7,1,1,7,4,12,59,0,2,59,1,1,60,0,1,60,2,1,
/* out0014_em-eta14-phi0*/	7,2,3,1,3,2,16,3,3,9,6,1,4,6,4,16,7,1,15,59,0,6,
/* out0015_em-eta15-phi0*/	5,2,2,3,2,3,6,3,3,7,3,4,4,59,0,3,
/* out0016_em-eta16-phi0*/	4,2,2,12,3,0,13,3,4,12,58,0,1,
/* out0017_em-eta17-phi0*/	5,2,1,3,2,2,1,3,0,3,3,1,7,58,0,4,
/* out0018_em-eta18-phi0*/	4,0,4,7,1,1,14,2,4,16,3,1,6,
/* out0019_em-eta19-phi0*/	6,0,2,15,0,3,15,0,4,1,0,5,1,1,0,12,1,1,2,
/* out0020_em-eta0-phi1*/	1,149,1,6,
/* out0021_em-eta1-phi1*/	2,148,3,3,149,1,10,
/* out0022_em-eta2-phi1*/	2,148,2,5,148,3,13,
/* out0023_em-eta3-phi1*/	8,60,1,12,60,2,9,70,0,4,70,1,2,71,1,3,71,2,12,147,3,6,148,2,11,
/* out0024_em-eta4-phi1*/	8,59,0,1,59,1,14,59,2,4,60,2,5,69,0,1,70,0,10,147,2,7,147,3,10,
/* out0025_em-eta5-phi1*/	6,58,0,1,58,1,12,59,2,11,69,0,6,146,3,8,147,2,9,
/* out0026_em-eta6-phi1*/	10,57,1,2,58,0,4,58,1,3,58,2,15,68,0,1,57,1,1,63,1,1,63,2,2,146,2,16,146,3,8,
/* out0027_em-eta7-phi1*/	8,57,0,6,57,1,11,57,2,3,57,0,13,57,1,1,62,1,4,63,1,9,63,2,1,
/* out0028_em-eta8-phi1*/	10,49,1,3,49,2,3,56,0,1,56,1,5,57,0,3,57,2,8,56,0,4,57,0,1,62,1,6,62,2,10,
/* out0029_em-eta9-phi1*/	6,56,0,9,56,1,3,56,2,2,56,0,4,61,1,12,62,2,2,
/* out0030_em-eta10-phi1*/	9,19,2,11,19,3,2,48,1,1,48,2,1,56,0,3,56,2,4,55,0,1,61,1,1,61,2,13,
/* out0031_em-eta11-phi1*/	8,18,5,3,19,0,4,19,2,5,19,3,1,19,4,9,19,5,14,48,2,1,60,1,11,
/* out0032_em-eta12-phi1*/	7,6,0,5,6,3,2,18,4,11,18,5,11,19,0,3,60,0,2,60,2,8,
/* out0033_em-eta13-phi1*/	7,6,0,10,6,1,3,17,2,10,17,5,3,18,4,1,59,1,6,60,2,2,
/* out0034_em-eta14-phi1*/	7,2,3,1,6,1,2,16,5,8,17,5,12,59,0,3,59,1,2,59,2,1,
/* out0035_em-eta15-phi1*/	6,2,0,3,2,3,7,16,4,3,16,5,5,59,0,2,59,2,5,
/* out0036_em-eta16-phi1*/	5,2,0,11,2,1,3,2,3,1,58,0,2,58,1,4,
/* out0037_em-eta17-phi1*/	6,2,0,1,2,1,9,3,1,2,5,2,1,5,5,3,58,0,5,
/* out0038_em-eta18-phi1*/	5,0,4,5,2,1,1,3,1,1,4,5,3,5,5,2,
/* out0039_em-eta19-phi1*/	7,0,2,1,0,3,1,0,4,3,0,5,11,1,0,4,1,3,16,1,5,16,
/* out0040_em-eta0-phi2*/	1,153,0,6,
/* out0041_em-eta1-phi2*/	2,152,0,3,153,0,10,
/* out0042_em-eta2-phi2*/	4,71,2,1,82,1,2,152,0,13,152,1,5,
/* out0043_em-eta3-phi2*/	8,70,1,13,71,1,13,71,2,3,82,0,16,82,1,2,82,2,1,151,0,6,152,1,11,
/* out0044_em-eta4-phi2*/	7,69,1,9,70,0,2,70,1,1,70,2,16,81,0,7,151,0,10,151,1,7,
/* out0045_em-eta5-phi2*/	6,68,1,1,69,0,9,69,1,6,69,2,13,150,0,8,151,1,9,
/* out0046_em-eta6-phi2*/	7,58,2,1,68,0,11,68,1,9,68,2,2,57,1,4,150,0,8,150,1,16,
/* out0047_em-eta7-phi2*/	10,57,1,3,57,2,3,67,0,2,67,1,3,68,0,4,68,2,4,50,0,1,57,0,2,57,1,10,57,2,12,
/* out0048_em-eta8-phi2*/	8,56,1,3,57,2,2,67,0,11,50,0,1,56,0,3,56,1,13,56,2,1,57,2,4,
/* out0049_em-eta9-phi2*/	7,56,1,5,56,2,6,66,0,1,67,0,1,55,1,2,56,0,5,56,2,10,
/* out0050_em-eta10-phi2*/	7,18,3,9,19,3,11,56,2,4,66,0,3,55,0,9,55,1,5,61,2,1,
/* out0051_em-eta11-phi2*/	12,18,0,2,18,1,3,18,2,15,18,3,7,19,0,3,19,3,2,19,4,7,54,1,1,55,0,6,55,2,3,60,1,3,60,2,1,
/* out0052_em-eta12-phi2*/	8,17,3,2,18,1,4,18,2,1,18,4,4,19,0,6,19,1,15,54,0,6,60,2,4,
/* out0053_em-eta13-phi2*/	7,16,2,1,17,2,6,17,3,12,17,4,7,17,5,1,54,0,4,59,1,4,
/* out0054_em-eta14-phi2*/	6,16,2,2,16,5,1,17,0,11,17,4,9,59,1,3,59,2,4,
/* out0055_em-eta15-phi2*/	6,16,4,11,16,5,2,17,0,2,17,1,3,53,0,1,59,2,5,
/* out0056_em-eta16-phi2*/	4,2,0,1,5,2,12,16,4,2,58,1,7,
/* out0057_em-eta17-phi2*/	5,5,2,2,5,4,2,5,5,9,58,0,3,58,1,1,
/* out0058_em-eta18-phi2*/	4,4,5,7,5,0,1,5,4,1,5,5,2,
/* out0059_em-eta19-phi2*/	3,0,5,4,4,4,4,4,5,4,
/* out0060_em-eta0-phi3*/	1,153,1,6,
/* out0061_em-eta1-phi3*/	2,152,3,3,153,1,10,
/* out0062_em-eta2-phi3*/	3,82,1,4,152,2,5,152,3,13,
/* out0063_em-eta3-phi3*/	7,81,1,5,82,1,8,82,2,15,124,0,11,124,1,3,151,3,6,152,2,11,
/* out0064_em-eta4-phi3*/	5,81,0,9,81,1,11,81,2,14,151,2,7,151,3,10,
/* out0065_em-eta5-phi3*/	8,69,1,1,69,2,3,80,0,13,80,1,10,80,2,2,81,2,1,150,3,8,151,2,9,
/* out0066_em-eta6-phi3*/	9,68,1,6,68,2,6,79,0,4,79,1,2,80,0,3,80,2,3,52,1,2,150,2,16,150,3,8,
/* out0067_em-eta7-phi3*/	8,67,1,10,68,2,4,79,0,6,50,0,7,50,1,13,50,2,2,52,0,1,52,1,1,
/* out0068_em-eta8-phi3*/	9,67,0,2,67,1,3,67,2,12,49,0,1,49,1,3,50,0,7,50,2,7,56,1,3,56,2,1,
/* out0069_em-eta9-phi3*/	7,66,0,3,66,1,9,67,2,2,49,0,12,49,1,1,55,1,2,56,2,4,
/* out0070_em-eta10-phi3*/	5,66,0,8,66,2,3,49,0,1,55,1,7,55,2,6,
/* out0071_em-eta11-phi3*/	9,18,0,14,18,1,2,21,2,13,21,5,2,66,0,1,66,2,1,48,0,1,54,1,4,55,2,7,
/* out0072_em-eta12-phi3*/	9,16,3,1,17,3,1,18,1,7,19,1,1,20,5,8,21,5,14,54,0,3,54,1,7,54,2,1,
/* out0073_em-eta13-phi3*/	8,16,0,4,16,2,3,16,3,15,17,3,1,20,4,1,20,5,3,54,0,3,54,2,5,
/* out0074_em-eta14-phi3*/	8,16,0,3,16,1,7,16,2,10,17,0,2,53,0,3,53,1,3,54,2,1,59,2,1,
/* out0075_em-eta15-phi3*/	5,5,3,2,16,1,3,17,0,1,17,1,13,53,0,6,
/* out0076_em-eta16-phi3*/	5,5,2,1,5,3,12,5,4,2,53,0,3,58,1,3,
/* out0077_em-eta17-phi3*/	5,4,2,2,5,0,1,5,4,11,58,0,1,58,1,1,
/* out0078_em-eta18-phi3*/	2,4,5,1,5,0,10,
/* out0079_em-eta19-phi3*/	3,4,4,7,4,5,1,5,1,1,
/* out0080_em-eta0-phi4*/	1,157,0,6,
/* out0081_em-eta1-phi4*/	2,156,0,3,157,0,10,
/* out0082_em-eta2-phi4*/	5,126,0,3,126,1,13,126,2,1,156,0,13,156,1,5,
/* out0083_em-eta3-phi4*/	9,124,0,4,124,1,13,124,2,14,125,1,1,125,2,6,126,0,13,126,2,5,155,0,6,156,1,11,
/* out0084_em-eta4-phi4*/	9,81,2,1,123,0,13,123,1,14,123,2,5,124,0,1,124,2,2,125,1,1,155,0,10,155,1,7,
/* out0085_em-eta5-phi4*/	8,80,1,6,80,2,8,122,0,6,122,1,3,123,0,3,123,2,4,154,0,8,155,1,9,
/* out0086_em-eta6-phi4*/	8,79,0,1,79,1,14,79,2,2,80,2,3,122,0,5,52,1,10,154,0,8,154,1,16,
/* out0087_em-eta7-phi4*/	10,78,1,3,79,0,5,79,2,11,50,1,3,50,2,3,51,1,3,51,2,4,52,0,15,52,1,2,52,2,11,
/* out0088_em-eta8-phi4*/	6,67,2,2,78,0,11,78,1,3,49,1,8,50,2,4,51,1,10,
/* out0089_em-eta9-phi4*/	6,66,1,7,66,2,2,78,0,5,49,0,2,49,1,4,49,2,12,
/* out0090_em-eta10-phi4*/	6,21,3,1,66,2,10,88,1,1,48,0,3,48,1,8,49,2,3,
/* out0091_em-eta11-phi4*/	8,20,2,4,20,3,6,21,2,3,21,3,15,21,4,8,48,0,11,48,2,1,54,1,1,
/* out0092_em-eta12-phi4*/	10,20,2,4,20,5,3,21,0,15,21,1,1,21,4,8,44,1,1,48,0,1,48,2,1,54,1,3,54,2,4,
/* out0093_em-eta13-phi4*/	9,16,0,4,20,4,14,20,5,2,21,1,2,28,5,1,29,5,3,44,1,2,53,1,1,54,2,5,
/* out0094_em-eta14-phi4*/	5,16,0,5,16,1,3,28,4,1,28,5,10,53,1,7,
/* out0095_em-eta15-phi4*/	7,4,3,1,5,3,1,16,1,3,28,4,11,53,0,2,53,1,1,53,2,3,
/* out0096_em-eta16-phi4*/	6,4,2,1,4,3,13,5,3,1,28,4,1,53,0,1,53,2,3,
/* out0097_em-eta17-phi4*/	3,4,1,1,4,2,10,4,3,2,
/* out0098_em-eta18-phi4*/	4,4,1,1,4,2,3,5,0,4,5,1,2,
/* out0099_em-eta19-phi4*/	2,4,4,5,5,1,8,
/* out0100_em-eta0-phi5*/	1,157,1,6,
/* out0101_em-eta1-phi5*/	2,156,3,3,157,1,10,
/* out0102_em-eta2-phi5*/	4,126,1,3,126,2,5,156,2,5,156,3,13,
/* out0103_em-eta3-phi5*/	6,125,0,16,125,1,7,125,2,10,126,2,5,155,3,6,156,2,11,
/* out0104_em-eta4-phi5*/	7,123,1,2,123,2,6,125,1,7,134,0,11,134,1,8,155,2,7,155,3,10,
/* out0105_em-eta5-phi5*/	7,122,0,2,122,1,13,122,2,7,123,2,1,134,0,5,154,3,8,155,2,9,
/* out0106_em-eta6-phi5*/	11,79,2,1,122,0,3,122,2,9,132,1,2,132,2,7,52,1,1,52,2,1,70,0,3,70,2,3,154,2,16,154,3,8,
/* out0107_em-eta7-phi5*/	9,78,1,4,79,2,2,132,1,13,51,0,2,51,2,12,52,2,4,70,0,2,70,1,8,70,2,13,
/* out0108_em-eta8-phi5*/	5,78,1,6,78,2,10,51,0,14,51,1,3,68,2,4,
/* out0109_em-eta9-phi5*/	6,78,2,6,88,1,1,88,2,7,49,2,1,68,1,12,68,2,4,
/* out0110_em-eta10-phi5*/	5,88,1,11,88,2,1,48,1,8,48,2,2,68,1,4,
/* out0111_em-eta11-phi5*/	6,20,0,13,20,2,2,20,3,10,88,1,3,44,2,1,48,2,11,
/* out0112_em-eta12-phi5*/	8,20,0,3,20,1,16,20,2,6,21,0,1,21,1,5,44,1,2,44,2,7,48,2,1,
/* out0113_em-eta13-phi5*/	5,20,4,1,21,1,8,29,2,7,29,5,9,44,1,9,
/* out0114_em-eta14-phi5*/	7,28,5,4,29,0,7,29,4,7,29,5,4,44,1,2,53,1,4,53,2,1,
/* out0115_em-eta15-phi5*/	5,28,4,2,28,5,1,29,0,8,29,1,7,53,2,6,
/* out0116_em-eta16-phi5*/	4,4,0,6,28,4,1,29,1,8,53,2,3,
/* out0117_em-eta17-phi5*/	2,4,0,10,4,1,3,
/* out0118_em-eta18-phi5*/	1,4,1,10,
/* out0119_em-eta19-phi5*/	2,4,1,1,5,1,5,
/* out0120_em-eta0-phi6*/	1,161,0,6,
/* out0121_em-eta1-phi6*/	2,160,0,3,161,0,10,
/* out0122_em-eta2-phi6*/	4,138,0,3,138,2,13,160,0,13,160,1,5,
/* out0123_em-eta3-phi6*/	7,136,0,15,136,1,6,136,2,5,138,1,4,138,2,3,159,0,6,160,1,11,
/* out0124_em-eta4-phi6*/	8,134,1,8,134,2,11,135,1,6,135,2,2,136,1,4,136,2,11,159,0,10,159,1,7,
/* out0125_em-eta5-phi6*/	7,133,0,2,133,1,7,133,2,13,134,2,5,135,1,1,158,0,8,159,1,9,
/* out0126_em-eta6-phi6*/	9,90,1,1,132,0,2,132,2,8,133,0,3,133,1,9,70,0,4,71,1,2,158,0,8,158,1,16,
/* out0127_em-eta7-phi6*/	11,89,2,4,90,1,2,132,0,14,132,1,1,132,2,1,69,1,2,69,2,12,70,0,7,70,1,8,71,0,2,71,1,3,
/* out0128_em-eta8-phi6*/	5,89,1,10,89,2,6,68,2,4,69,0,3,69,1,14,
/* out0129_em-eta9-phi6*/	6,88,0,1,88,2,7,89,1,6,46,1,1,68,0,12,68,2,4,
/* out0130_em-eta10-phi6*/	5,88,0,10,88,2,1,45,1,2,45,2,8,68,0,4,
/* out0131_em-eta11-phi6*/	7,30,5,5,31,2,3,31,4,2,31,5,15,88,0,3,44,2,1,45,1,11,
/* out0132_em-eta12-phi6*/	7,30,4,10,30,5,11,31,0,7,31,1,2,44,0,2,44,2,7,45,1,1,
/* out0133_em-eta13-phi6*/	5,29,2,9,29,3,8,30,4,6,31,1,4,44,0,8,
/* out0134_em-eta14-phi6*/	7,28,2,7,28,3,2,29,3,4,29,4,9,39,1,1,39,2,4,44,0,2,
/* out0135_em-eta15-phi6*/	6,28,0,1,28,1,7,28,2,9,28,3,1,29,0,1,39,1,6,
/* out0136_em-eta16-phi6*/	4,28,1,9,29,1,1,37,5,6,39,1,3,
/* out0137_em-eta17-phi6*/	2,36,5,11,37,5,2,
/* out0138_em-eta18-phi6*/	2,36,4,7,36,5,3,
/* out0139_em-eta19-phi6*/	1,36,4,5,
/* out0140_em-eta0-phi7*/	1,161,1,6,
/* out0141_em-eta1-phi7*/	2,160,3,3,161,1,10,
/* out0142_em-eta2-phi7*/	4,138,0,13,138,1,1,160,2,5,160,3,13,
/* out0143_em-eta3-phi7*/	8,136,0,1,136,1,6,137,0,4,137,1,14,137,2,13,138,1,11,159,3,6,160,2,11,
/* out0144_em-eta4-phi7*/	8,92,1,1,135,0,13,135,1,5,135,2,14,137,0,1,137,1,2,159,2,7,159,3,10,
/* out0145_em-eta5-phi7*/	8,91,1,8,91,2,6,133,0,6,133,2,3,135,0,3,135,1,4,158,3,8,159,2,9,
/* out0146_em-eta6-phi7*/	9,90,0,1,90,1,2,90,2,14,91,1,3,133,0,5,71,1,8,71,2,3,158,2,16,158,3,8,
/* out0147_em-eta7-phi7*/	10,89,2,3,90,0,5,90,1,11,47,1,3,47,2,3,69,0,3,69,2,4,71,0,14,71,1,3,71,2,10,
/* out0148_em-eta8-phi7*/	6,89,0,11,89,2,3,101,1,2,46,2,8,47,1,4,69,0,10,
/* out0149_em-eta9-phi7*/	6,89,0,5,100,1,2,100,2,7,46,0,2,46,1,12,46,2,4,
/* out0150_em-eta10-phi7*/	6,31,2,1,88,0,2,100,1,10,45,0,3,45,2,8,46,1,3,
/* out0151_em-eta11-phi7*/	9,30,2,1,30,3,1,31,2,12,31,3,11,31,4,10,31,5,1,40,2,1,45,0,11,45,1,1,
/* out0152_em-eta12-phi7*/	10,30,1,4,30,2,15,31,0,9,31,1,1,31,4,4,40,1,4,40,2,3,44,0,2,45,0,1,45,1,1,
/* out0153_em-eta13-phi7*/	9,28,3,1,29,3,3,30,1,9,31,1,9,38,5,1,39,5,3,39,2,1,40,1,5,44,0,2,
/* out0154_em-eta14-phi7*/	6,28,0,1,28,3,12,29,3,1,38,4,1,38,5,7,39,2,7,
/* out0155_em-eta15-phi7*/	6,28,0,13,37,2,2,38,4,3,39,0,2,39,1,3,39,2,1,
/* out0156_em-eta16-phi7*/	6,28,0,1,37,2,7,37,4,1,37,5,6,39,0,1,39,1,3,
/* out0157_em-eta17-phi7*/	4,36,5,1,37,0,5,37,4,6,37,5,2,
/* out0158_em-eta18-phi7*/	4,36,4,1,36,5,1,37,0,7,37,1,2,
/* out0159_em-eta19-phi7*/	2,36,4,3,37,1,7,
/* out0160_em-eta0-phi8*/	1,165,0,6,
/* out0161_em-eta1-phi8*/	2,164,0,3,165,0,10,
/* out0162_em-eta2-phi8*/	3,93,2,4,164,0,13,164,1,5,
/* out0163_em-eta3-phi8*/	7,92,2,5,93,1,15,93,2,8,137,0,11,137,2,3,163,0,6,164,1,11,
/* out0164_em-eta4-phi8*/	5,92,0,9,92,1,14,92,2,11,163,0,10,163,1,7,
/* out0165_em-eta5-phi8*/	8,91,0,13,91,1,2,91,2,10,92,1,1,103,1,3,103,2,1,162,0,8,163,1,9,
/* out0166_em-eta6-phi8*/	9,90,0,4,90,2,2,91,0,3,91,1,3,102,1,6,102,2,6,71,2,2,162,0,8,162,1,16,
/* out0167_em-eta7-phi8*/	7,90,0,6,101,2,10,102,1,4,47,0,7,47,1,2,47,2,13,71,2,1,
/* out0168_em-eta8-phi8*/	9,101,0,2,101,1,12,101,2,3,42,1,1,42,2,3,46,0,1,46,2,3,47,0,7,47,1,7,
/* out0169_em-eta9-phi8*/	7,100,0,3,100,2,9,101,1,2,41,2,2,42,1,4,46,0,12,46,2,1,
/* out0170_em-eta10-phi8*/	5,100,0,8,100,1,3,41,1,6,41,2,7,46,0,1,
/* out0171_em-eta11-phi8*/	9,30,3,9,31,3,5,40,5,10,41,5,7,100,0,1,100,1,1,40,2,4,41,1,7,45,0,1,
/* out0172_em-eta12-phi8*/	9,30,0,14,30,1,1,30,3,6,39,2,2,40,4,7,40,5,1,40,0,3,40,1,1,40,2,7,
/* out0173_em-eta13-phi8*/	7,30,0,2,30,1,2,39,2,8,39,4,3,39,5,12,40,0,3,40,1,5,
/* out0174_em-eta14-phi8*/	9,38,4,1,38,5,8,39,0,9,39,4,3,39,5,1,34,1,1,39,0,3,39,2,3,40,1,1,
/* out0175_em-eta15-phi8*/	5,37,2,2,38,4,11,39,0,1,39,1,5,39,0,6,
/* out0176_em-eta16-phi8*/	5,37,2,5,37,3,9,37,4,2,33,1,3,39,0,3,
/* out0177_em-eta17-phi8*/	3,36,2,5,37,4,7,33,1,2,
/* out0178_em-eta18-phi8*/	4,36,1,1,36,2,6,37,0,4,37,1,2,
/* out0179_em-eta19-phi8*/	2,36,1,5,37,1,5,
/* out0180_em-eta0-phi9*/	1,165,1,6,
/* out0181_em-eta1-phi9*/	2,164,3,3,165,1,10,
/* out0182_em-eta2-phi9*/	4,93,2,2,105,0,1,164,2,5,164,3,13,
/* out0183_em-eta3-phi9*/	8,93,0,16,93,1,1,93,2,2,104,2,13,105,0,3,105,1,13,163,3,6,164,2,11,
/* out0184_em-eta4-phi9*/	7,92,0,7,103,2,9,104,0,2,104,1,16,104,2,1,163,2,7,163,3,10,
/* out0185_em-eta5-phi9*/	6,102,2,1,103,0,9,103,1,13,103,2,6,162,3,8,163,2,9,
/* out0186_em-eta6-phi9*/	7,102,0,11,102,1,2,102,2,9,114,1,1,43,2,4,162,2,16,162,3,8,
/* out0187_em-eta7-phi9*/	10,101,0,2,101,2,3,102,0,4,102,1,4,113,1,3,113,2,3,43,0,2,43,1,12,43,2,10,47,0,1,
/* out0188_em-eta8-phi9*/	8,101,0,11,112,2,3,113,1,2,42,0,3,42,1,1,42,2,13,43,1,4,47,0,1,
/* out0189_em-eta9-phi9*/	7,100,0,1,101,0,1,112,1,6,112,2,5,41,2,2,42,0,5,42,1,10,
/* out0190_em-eta10-phi9*/	8,41,2,16,41,3,3,41,5,1,100,0,3,112,1,4,36,1,1,41,0,9,41,2,5,
/* out0191_em-eta11-phi9*/	11,40,2,2,40,5,3,41,0,9,41,3,1,41,4,14,41,5,8,35,1,1,35,2,3,40,2,1,41,0,6,41,1,3,
/* out0192_em-eta12-phi9*/	7,39,2,2,40,4,9,40,5,2,41,0,7,41,1,12,35,1,4,40,0,6,
/* out0193_em-eta13-phi9*/	7,38,2,1,38,3,1,39,2,4,39,3,14,39,4,7,34,2,4,40,0,4,
/* out0194_em-eta14-phi9*/	6,38,1,1,38,2,13,39,0,4,39,4,3,34,1,4,34,2,3,
/* out0195_em-eta15-phi9*/	6,38,1,7,38,2,1,39,0,2,39,1,9,34,1,5,39,0,1,
/* out0196_em-eta16-phi9*/	5,36,3,6,37,3,7,39,1,2,33,1,4,33,2,3,
/* out0197_em-eta17-phi9*/	4,36,0,1,36,2,3,36,3,9,33,1,4,
/* out0198_em-eta18-phi9*/	3,36,0,5,36,1,4,36,2,2,
/* out0199_em-eta19-phi9*/	3,8,3,3,36,0,1,36,1,6,
/* out0200_em-eta0-phi10*/	1,169,0,6,
/* out0201_em-eta1-phi10*/	2,168,0,3,169,0,10,
/* out0202_em-eta2-phi10*/	2,168,0,13,168,1,5,
/* out0203_em-eta3-phi10*/	8,104,0,4,104,2,2,105,0,12,105,1,3,116,1,9,116,2,12,167,0,6,168,1,11,
/* out0204_em-eta4-phi10*/	8,103,0,1,104,0,10,115,0,1,115,1,4,115,2,14,116,1,5,167,0,10,167,1,7,
/* out0205_em-eta5-phi10*/	6,103,0,6,114,0,1,114,2,12,115,1,11,166,0,8,167,1,9,
/* out0206_em-eta6-phi10*/	10,102,0,1,113,2,2,114,0,4,114,1,15,114,2,3,38,0,2,38,1,1,43,2,1,166,0,8,166,1,16,
/* out0207_em-eta7-phi10*/	8,113,0,6,113,1,3,113,2,11,37,2,4,38,0,1,38,1,9,43,0,13,43,2,1,
/* out0208_em-eta8-phi10*/	8,112,0,1,112,2,5,113,0,3,113,1,8,37,1,10,37,2,6,42,0,4,43,0,1,
/* out0209_em-eta9-phi10*/	6,112,0,9,112,1,2,112,2,3,36,2,12,37,1,2,42,0,4,
/* out0210_em-eta10-phi10*/	8,40,3,3,41,3,10,52,0,2,112,0,3,112,1,4,36,1,13,36,2,1,41,0,1,
/* out0211_em-eta11-phi10*/	7,40,0,8,40,1,1,40,2,11,40,3,13,41,3,2,41,4,2,35,2,11,
/* out0212_em-eta12-phi10*/	7,15,5,5,40,0,4,40,1,15,40,2,3,41,1,3,35,0,2,35,1,8,
/* out0213_em-eta13-phi10*/	8,14,4,1,14,5,9,15,5,2,38,3,11,39,3,2,41,1,1,34,2,6,35,1,2,
/* out0214_em-eta14-phi10*/	8,14,4,1,38,0,14,38,1,2,38,2,1,38,3,4,34,0,3,34,1,1,34,2,2,
/* out0215_em-eta15-phi10*/	6,13,2,3,13,5,7,38,0,2,38,1,6,34,0,2,34,1,5,
/* out0216_em-eta16-phi10*/	3,12,5,10,13,5,5,33,2,6,
/* out0217_em-eta17-phi10*/	6,12,4,5,12,5,3,36,0,3,36,3,1,33,1,2,33,2,2,
/* out0218_em-eta18-phi10*/	3,8,0,4,12,4,1,36,0,6,
/* out0219_em-eta19-phi10*/	6,8,0,3,8,2,1,8,3,11,8,5,1,9,3,16,9,5,16,
/* out0220_em-eta0-phi11*/	1,169,1,6,
/* out0221_em-eta1-phi11*/	2,168,3,3,169,1,10,
/* out0222_em-eta2-phi11*/	2,168,2,5,168,3,13,
/* out0223_em-eta3-phi11*/	4,116,0,14,116,2,4,167,3,6,168,2,11,
/* out0224_em-eta4-phi11*/	7,55,1,1,115,0,10,115,2,2,116,0,2,116,1,2,167,2,7,167,3,10,
/* out0225_em-eta5-phi11*/	9,55,0,15,55,1,3,55,2,1,114,0,3,114,2,1,115,0,5,115,1,1,166,3,8,167,2,9,
/* out0226_em-eta6-phi11*/	8,54,0,8,54,1,4,55,0,1,55,2,2,114,0,8,38,0,1,166,2,16,166,3,8,
/* out0227_em-eta7-phi11*/	9,53,1,2,54,0,8,54,2,4,113,0,6,32,0,6,37,0,1,37,2,4,38,0,12,38,1,6,
/* out0228_em-eta8-phi11*/	8,53,0,12,53,1,2,113,0,1,31,0,2,32,0,1,37,0,14,37,1,2,37,2,2,
/* out0229_em-eta9-phi11*/	10,52,0,1,52,1,2,53,0,4,53,2,4,112,0,3,31,0,6,36,0,6,36,2,3,37,0,1,37,1,2,
/* out0230_em-eta10-phi11*/	5,52,0,9,52,1,2,30,0,3,36,0,10,36,1,2,
/* out0231_em-eta11-phi11*/	7,15,2,3,40,0,3,52,0,4,52,2,4,30,0,5,35,0,5,35,2,2,
/* out0232_em-eta12-phi11*/	7,15,2,13,15,3,3,15,4,7,15,5,7,40,0,1,29,0,2,35,0,8,
/* out0233_em-eta13-phi11*/	11,14,4,1,14,5,7,15,0,12,15,1,1,15,4,4,15,5,2,29,0,5,34,0,2,34,2,1,35,0,1,35,1,1,
/* out0234_em-eta14-phi11*/	5,13,2,6,14,4,13,15,1,3,29,0,1,34,0,6,
/* out0235_em-eta15-phi11*/	6,13,2,7,13,3,3,13,4,5,13,5,3,28,0,3,34,0,3,
/* out0236_em-eta16-phi11*/	6,12,5,1,13,0,8,13,4,6,13,5,1,28,0,4,33,2,2,
/* out0237_em-eta17-phi11*/	7,12,4,5,12,5,2,13,0,3,13,1,3,28,0,1,33,1,1,33,2,3,
/* out0238_em-eta18-phi11*/	4,8,0,7,8,1,2,12,4,5,13,1,1,
/* out0239_em-eta19-phi11*/	6,8,0,2,8,1,2,8,2,11,8,3,2,8,5,13,9,0,4,
/* out0240_em-eta0-phi12*/	1,173,0,6,
/* out0241_em-eta1-phi12*/	2,172,0,3,173,0,10,
/* out0242_em-eta2-phi12*/	2,172,0,13,172,1,5,
/* out0243_em-eta3-phi12*/	4,65,0,14,65,1,4,171,0,6,172,1,11,
/* out0244_em-eta4-phi12*/	7,55,1,1,64,0,10,64,1,2,65,0,2,65,2,2,171,0,10,171,1,7,
/* out0245_em-eta5-phi12*/	8,55,1,11,55,2,9,63,0,3,63,1,1,64,0,5,64,2,1,170,0,8,171,1,9,
/* out0246_em-eta6-phi12*/	6,54,1,12,55,2,4,63,0,8,32,1,1,170,0,8,170,1,16,
/* out0247_em-eta7-phi12*/	6,53,1,2,54,2,12,62,0,6,32,0,7,32,1,13,32,2,5,
/* out0248_em-eta8-phi12*/	7,53,1,10,53,2,5,62,0,1,31,0,2,31,1,10,32,0,2,32,2,8,
/* out0249_em-eta9-phi12*/	6,52,1,3,53,2,7,61,0,3,31,0,6,31,1,2,31,2,9,
/* out0250_em-eta10-phi12*/	5,52,1,8,52,2,3,30,0,3,30,1,9,31,2,2,
/* out0251_em-eta11-phi12*/	7,15,3,3,26,5,1,27,5,2,52,2,8,30,0,5,30,1,1,30,2,7,
/* out0252_em-eta12-phi12*/	8,14,2,4,14,3,13,15,3,10,15,4,4,26,5,1,29,0,2,29,1,6,30,2,2,
/* out0253_em-eta13-phi12*/	10,14,0,1,14,1,7,14,2,12,14,3,1,15,0,4,15,1,1,15,4,1,29,0,5,29,1,1,29,2,3,
/* out0254_em-eta14-phi12*/	7,12,3,1,13,3,6,14,1,4,15,1,11,28,1,2,29,0,1,29,2,4,
/* out0255_em-eta15-phi12*/	6,12,2,3,12,3,6,13,3,7,13,4,4,28,0,3,28,1,3,
/* out0256_em-eta16-phi12*/	5,12,2,12,13,0,2,13,4,1,28,0,4,28,2,1,
/* out0257_em-eta17-phi12*/	6,12,1,3,12,2,1,13,0,3,13,1,6,28,0,1,28,2,3,
/* out0258_em-eta18-phi12*/	3,8,1,10,9,1,1,13,1,5,
/* out0259_em-eta19-phi12*/	6,8,1,1,8,2,4,8,4,7,8,5,2,9,0,12,9,1,4,
/* out0260_em-eta0-phi13*/	1,173,1,6,
/* out0261_em-eta1-phi13*/	2,172,3,3,173,1,10,
/* out0262_em-eta2-phi13*/	2,172,2,5,172,3,13,
/* out0263_em-eta3-phi13*/	8,65,1,12,65,2,9,76,0,4,76,1,2,77,0,12,77,2,3,171,3,6,172,2,11,
/* out0264_em-eta4-phi13*/	8,64,0,1,64,1,14,64,2,4,65,2,5,75,0,1,76,0,10,171,2,7,171,3,10,
/* out0265_em-eta5-phi13*/	6,63,0,1,63,1,12,64,2,11,75,0,6,170,3,8,171,2,9,
/* out0266_em-eta6-phi13*/	8,62,1,2,63,0,4,63,1,3,63,2,15,74,0,1,27,0,5,170,2,16,170,3,8,
/* out0267_em-eta7-phi13*/	9,62,0,6,62,1,11,62,2,3,26,0,3,26,1,6,27,0,10,27,2,9,32,1,2,32,2,2,
/* out0268_em-eta8-phi13*/	9,61,0,1,61,1,5,62,0,3,62,2,8,26,0,13,26,1,2,26,2,4,31,1,2,32,2,1,
/* out0269_em-eta9-phi13*/	8,61,0,9,61,1,3,61,2,2,25,0,7,25,1,3,26,2,1,31,1,2,31,2,5,
/* out0270_em-eta10-phi13*/	9,27,2,11,27,3,2,52,1,1,52,2,1,61,0,3,61,2,4,25,0,8,25,2,1,30,1,6,
/* out0271_em-eta11-phi13*/	8,26,5,3,27,0,4,27,2,5,27,3,1,27,4,9,27,5,14,24,0,5,30,2,7,
/* out0272_em-eta12-phi13*/	7,14,0,5,14,3,2,26,4,11,26,5,11,27,0,3,24,0,4,29,1,6,
/* out0273_em-eta13-phi13*/	7,14,0,10,14,1,3,23,2,10,23,5,3,26,4,1,29,1,3,29,2,6,
/* out0274_em-eta14-phi13*/	8,12,3,1,14,1,2,22,5,8,23,4,1,23,5,12,23,0,1,28,1,2,29,2,3,
/* out0275_em-eta15-phi13*/	5,12,0,3,12,3,7,22,4,3,22,5,5,28,1,6,
/* out0276_em-eta16-phi13*/	5,12,0,11,12,1,3,12,3,1,28,1,1,28,2,5,
/* out0277_em-eta17-phi13*/	5,11,2,1,11,5,3,12,0,1,12,1,9,28,2,3,
/* out0278_em-eta18-phi13*/	6,8,1,1,9,1,5,10,5,3,11,5,2,12,1,1,13,1,1,
/* out0279_em-eta19-phi13*/	2,8,4,6,9,1,6,
/* out0280_em-eta0-phi14*/	1,177,0,6,
/* out0281_em-eta1-phi14*/	2,176,0,3,177,0,10,
/* out0282_em-eta2-phi14*/	4,77,0,1,87,1,2,176,0,13,176,1,5,
/* out0283_em-eta3-phi14*/	8,76,1,13,77,0,3,77,2,13,87,0,16,87,1,2,87,2,1,175,0,6,176,1,11,
/* out0284_em-eta4-phi14*/	7,75,1,9,76,0,2,76,1,1,76,2,16,86,0,7,175,0,10,175,1,7,
/* out0285_em-eta5-phi14*/	6,74,1,1,75,0,9,75,1,6,75,2,14,174,0,8,175,1,9,
/* out0286_em-eta6-phi14*/	10,63,2,1,74,0,11,74,1,9,74,2,2,21,0,4,21,2,1,27,0,1,27,2,2,174,0,8,174,1,16,
/* out0287_em-eta7-phi14*/	11,62,1,3,62,2,3,73,0,2,73,1,3,74,0,4,74,2,4,21,0,4,21,1,3,21,2,15,26,1,5,27,2,5,
/* out0288_em-eta8-phi14*/	7,61,1,3,62,2,2,73,0,11,19,0,6,19,1,1,26,1,3,26,2,11,
/* out0289_em-eta9-phi14*/	7,61,1,5,61,2,6,72,0,1,73,0,1,19,0,2,25,1,13,25,2,2,
/* out0290_em-eta10-phi14*/	7,26,3,9,27,3,11,61,2,4,72,0,3,24,1,2,25,0,1,25,2,12,
/* out0291_em-eta11-phi14*/	10,26,0,2,26,1,3,26,2,15,26,3,7,27,0,3,27,3,2,27,4,7,24,0,3,24,1,9,24,2,1,
/* out0292_em-eta12-phi14*/	8,23,3,2,26,1,4,26,2,1,26,4,4,27,0,6,27,1,15,24,0,4,24,2,6,
/* out0293_em-eta13-phi14*/	7,22,2,1,23,2,6,23,3,12,23,4,7,23,5,1,23,0,4,23,1,4,
/* out0294_em-eta14-phi14*/	5,22,2,2,22,5,1,23,0,11,23,4,8,23,0,7,
/* out0295_em-eta15-phi14*/	6,22,4,11,22,5,2,23,0,2,23,1,3,23,0,3,28,1,2,
/* out0296_em-eta16-phi14*/	5,11,2,12,12,0,1,22,4,2,22,1,2,28,2,3,
/* out0297_em-eta17-phi14*/	6,11,2,2,11,4,2,11,5,9,22,0,1,22,1,2,28,2,1,
/* out0298_em-eta18-phi14*/	4,10,5,8,11,0,1,11,4,1,11,5,2,
/* out0299_em-eta19-phi14*/	3,8,4,3,10,4,4,10,5,3,
/* out0300_em-eta0-phi15*/	1,177,1,6,
/* out0301_em-eta1-phi15*/	2,176,3,3,177,1,10,
/* out0302_em-eta2-phi15*/	3,87,1,4,176,2,5,176,3,13,
/* out0303_em-eta3-phi15*/	7,86,1,5,87,1,8,87,2,15,130,0,11,130,1,3,175,3,6,176,2,11,
/* out0304_em-eta4-phi15*/	5,86,0,9,86,1,11,86,2,14,175,2,7,175,3,10,
/* out0305_em-eta5-phi15*/	8,75,1,1,75,2,2,85,0,13,85,1,10,85,2,2,86,2,1,174,3,8,175,2,9,
/* out0306_em-eta6-phi15*/	9,74,1,6,74,2,6,84,0,4,84,1,2,85,0,3,85,2,3,21,0,1,174,2,16,174,3,8,
/* out0307_em-eta7-phi15*/	7,73,1,10,74,2,4,84,0,6,19,1,1,20,1,6,21,0,7,21,1,13,
/* out0308_em-eta8-phi15*/	6,73,0,2,73,1,3,73,2,12,19,0,4,19,1,13,19,2,4,
/* out0309_em-eta9-phi15*/	8,72,0,3,72,1,9,73,2,2,17,0,1,17,1,5,19,0,4,19,2,7,25,2,1,
/* out0310_em-eta10-phi15*/	4,72,0,8,72,2,3,17,0,12,17,1,1,
/* out0311_em-eta11-phi15*/	11,25,2,13,25,5,2,26,0,14,26,1,2,72,0,1,72,2,1,16,0,1,17,0,3,17,2,1,24,1,5,24,2,3,
/* out0312_em-eta12-phi15*/	9,22,3,1,23,3,1,24,5,8,25,5,14,26,1,7,27,1,1,16,0,4,23,1,1,24,2,6,
/* out0313_em-eta13-phi15*/	7,22,0,4,22,2,3,22,3,15,23,3,1,24,4,1,24,5,3,23,1,8,
/* out0314_em-eta14-phi15*/	7,22,0,3,22,1,7,22,2,10,23,0,2,23,0,1,23,1,1,23,2,6,
/* out0315_em-eta15-phi15*/	6,11,3,2,22,1,3,23,0,1,23,1,13,22,1,2,23,2,4,
/* out0316_em-eta16-phi15*/	4,11,2,1,11,3,12,11,4,2,22,1,5,
/* out0317_em-eta17-phi15*/	5,10,2,2,11,0,1,11,4,11,22,0,4,22,1,1,
/* out0318_em-eta18-phi15*/	2,10,5,1,11,0,10,
/* out0319_em-eta19-phi15*/	3,10,4,7,10,5,1,11,1,1,
/* out0320_em-eta0-phi16*/	1,181,0,6,
/* out0321_em-eta1-phi16*/	2,180,0,3,181,0,10,
/* out0322_em-eta2-phi16*/	5,131,0,1,131,1,16,131,2,8,180,0,13,180,1,5,
/* out0323_em-eta3-phi16*/	8,129,1,1,129,2,6,130,0,4,130,1,13,130,2,14,131,0,11,179,0,6,180,1,11,
/* out0324_em-eta4-phi16*/	9,86,2,1,128,0,13,128,1,14,128,2,5,129,1,1,130,0,1,130,2,2,179,0,10,179,1,7,
/* out0325_em-eta5-phi16*/	8,85,1,6,85,2,8,127,0,6,127,1,3,128,0,3,128,2,4,178,0,8,179,1,9,
/* out0326_em-eta6-phi16*/	8,84,0,1,84,1,14,84,2,2,85,2,3,127,0,5,20,2,3,178,0,8,178,1,16,
/* out0327_em-eta7-phi16*/	6,83,1,3,84,0,5,84,2,11,20,0,7,20,1,7,20,2,12,
/* out0328_em-eta8-phi16*/	9,73,2,2,83,0,11,83,1,3,18,1,5,18,2,5,19,1,1,19,2,3,20,0,4,20,1,3,
/* out0329_em-eta9-phi16*/	6,72,1,7,72,2,2,83,0,5,17,1,6,18,1,10,19,2,2,
/* out0330_em-eta10-phi16*/	5,25,3,1,72,2,10,94,1,1,17,1,4,17,2,11,
/* out0331_em-eta11-phi16*/	8,24,2,4,24,3,6,25,2,3,25,3,15,25,4,8,16,0,1,16,1,8,17,2,4,
/* out0332_em-eta12-phi16*/	8,24,2,4,24,5,3,25,0,15,25,1,1,25,4,8,16,0,7,16,1,1,16,2,1,
/* out0333_em-eta13-phi16*/	11,22,0,4,24,4,14,24,5,2,25,1,2,32,5,1,33,5,3,11,1,1,16,0,3,16,2,2,23,1,2,23,2,1,
/* out0334_em-eta14-phi16*/	6,22,0,5,22,1,3,32,4,1,32,5,10,11,1,3,23,2,4,
/* out0335_em-eta15-phi16*/	8,10,3,1,11,3,1,22,1,3,32,4,11,11,1,1,22,1,2,22,2,2,23,2,1,
/* out0336_em-eta16-phi16*/	6,10,2,1,10,3,13,11,3,1,32,4,1,22,1,2,22,2,3,
/* out0337_em-eta17-phi16*/	5,10,1,1,10,2,10,10,3,2,22,0,6,22,2,1,
/* out0338_em-eta18-phi16*/	5,10,1,1,10,2,3,11,0,4,11,1,2,22,0,2,
/* out0339_em-eta19-phi16*/	2,10,4,5,11,1,8,
/* out0340_em-eta0-phi17*/	1,181,1,6,
/* out0341_em-eta1-phi17*/	2,180,3,3,181,1,10,
/* out0342_em-eta2-phi17*/	3,131,2,7,180,2,5,180,3,13,
/* out0343_em-eta3-phi17*/	7,129,0,16,129,1,7,129,2,10,131,0,4,131,2,1,179,3,6,180,2,11,
/* out0344_em-eta4-phi17*/	7,128,1,2,128,2,6,129,1,7,143,0,11,143,1,8,179,2,7,179,3,10,
/* out0345_em-eta5-phi17*/	7,127,0,2,127,1,13,127,2,7,128,2,1,143,0,5,178,3,8,179,2,9,
/* out0346_em-eta6-phi17*/	7,84,2,1,127,0,3,127,2,9,139,1,2,139,2,7,178,2,16,178,3,8,
/* out0347_em-eta7-phi17*/	7,83,1,4,84,2,2,139,1,13,20,0,4,20,2,1,67,0,10,67,1,7,
/* out0348_em-eta8-phi17*/	6,83,1,6,83,2,10,18,0,4,18,2,11,20,0,1,67,0,6,
/* out0349_em-eta9-phi17*/	6,83,2,6,94,1,1,94,2,7,18,0,12,18,1,1,64,2,4,
/* out0350_em-eta10-phi17*/	4,94,1,11,94,2,1,64,1,10,64,2,4,
/* out0351_em-eta11-phi17*/	7,24,0,13,24,2,2,24,3,10,94,1,3,16,1,6,16,2,1,64,1,6,
/* out0352_em-eta12-phi17*/	7,24,0,3,24,1,16,24,2,6,25,0,1,25,1,5,16,1,1,16,2,9,
/* out0353_em-eta13-phi17*/	6,24,4,1,25,1,8,33,2,7,33,5,9,11,2,5,16,2,3,
/* out0354_em-eta14-phi17*/	6,32,5,4,33,0,7,33,4,7,33,5,4,11,1,5,11,2,2,
/* out0355_em-eta15-phi17*/	6,32,4,2,32,5,1,33,0,8,33,1,7,11,1,6,22,2,1,
/* out0356_em-eta16-phi17*/	4,10,0,6,32,4,1,33,1,8,22,2,5,
/* out0357_em-eta17-phi17*/	4,10,0,10,10,1,3,22,0,1,22,2,4,
/* out0358_em-eta18-phi17*/	3,10,1,10,11,1,1,22,0,2,
/* out0359_em-eta19-phi17*/	2,10,1,1,11,1,4,
/* out0360_em-eta0-phi18*/	1,185,0,6,
/* out0361_em-eta1-phi18*/	2,184,0,3,185,0,10,
/* out0362_em-eta2-phi18*/	3,145,0,8,184,0,13,184,1,5,
/* out0363_em-eta3-phi18*/	7,144,0,16,144,1,11,144,2,5,145,0,1,145,2,10,183,0,6,184,1,11,
/* out0364_em-eta4-phi18*/	7,141,1,6,141,2,2,143,1,8,143,2,10,144,2,9,183,0,10,183,1,7,
/* out0365_em-eta5-phi18*/	7,140,0,2,140,1,7,140,2,13,141,1,1,143,2,6,182,0,8,183,1,9,
/* out0366_em-eta6-phi18*/	8,96,1,1,139,0,2,139,2,8,140,0,3,140,1,9,67,1,1,182,0,8,182,1,16,
/* out0367_em-eta7-phi18*/	9,95,2,4,96,1,2,139,0,14,139,1,1,139,2,1,66,1,4,66,2,1,67,1,8,67,2,10,
/* out0368_em-eta8-phi18*/	6,95,1,10,95,2,6,65,1,4,65,2,11,66,1,1,67,2,6,
/* out0369_em-eta9-phi18*/	6,94,0,1,94,2,7,95,1,6,64,2,4,65,0,1,65,1,12,
/* out0370_em-eta10-phi18*/	4,94,0,10,94,2,1,64,0,10,64,2,4,
/* out0371_em-eta11-phi18*/	8,34,5,5,35,2,3,35,4,2,35,5,15,94,0,3,12,1,1,12,2,6,64,0,6,
/* out0372_em-eta12-phi18*/	6,34,4,10,34,5,11,35,0,7,35,1,2,12,1,9,12,2,1,
/* out0373_em-eta13-phi18*/	6,33,2,9,33,3,8,34,4,6,35,1,4,11,2,6,12,1,3,
/* out0374_em-eta14-phi18*/	6,32,2,7,32,3,2,33,3,4,33,4,9,11,0,5,11,2,2,
/* out0375_em-eta15-phi18*/	6,32,0,1,32,1,7,32,2,9,32,3,1,33,0,1,11,0,5,
/* out0376_em-eta16-phi18*/	4,32,1,9,33,1,1,43,5,6,5,1,4,
/* out0377_em-eta17-phi18*/	3,42,5,11,43,5,2,5,1,4,
/* out0378_em-eta18-phi18*/	3,42,4,7,42,5,3,5,0,1,
/* out0379_em-eta19-phi18*/	1,42,4,5,
/* out0380_em-eta0-phi19*/	1,185,1,6,
/* out0381_em-eta1-phi19*/	2,184,3,3,185,1,10,
/* out0382_em-eta2-phi19*/	4,145,0,7,145,1,8,184,2,5,184,3,13,
/* out0383_em-eta3-phi19*/	9,142,0,4,142,1,14,142,2,13,144,1,5,144,2,1,145,1,8,145,2,6,183,3,6,184,2,11,
/* out0384_em-eta4-phi19*/	9,98,1,1,141,0,13,141,1,5,141,2,14,142,0,1,142,1,2,144,2,1,183,2,7,183,3,10,
/* out0385_em-eta5-phi19*/	8,97,1,8,97,2,6,140,0,6,140,2,3,141,0,3,141,1,4,182,3,8,183,2,9,
/* out0386_em-eta6-phi19*/	8,96,0,1,96,1,2,96,2,14,97,1,3,140,0,5,66,2,3,182,2,16,182,3,8,
/* out0387_em-eta7-phi19*/	6,95,2,3,96,0,5,96,1,11,66,0,7,66,1,7,66,2,12,
/* out0388_em-eta8-phi19*/	9,95,0,11,95,2,3,107,1,2,14,1,3,14,2,1,65,0,5,65,2,5,66,0,3,66,1,4,
/* out0389_em-eta9-phi19*/	6,95,0,5,106,1,2,106,2,7,13,2,6,14,1,2,65,0,10,
/* out0390_em-eta10-phi19*/	5,35,2,1,94,0,2,106,1,10,13,1,11,13,2,4,
/* out0391_em-eta11-phi19*/	9,34,2,1,34,3,1,35,2,12,35,3,11,35,4,10,35,5,1,12,0,1,12,2,8,13,1,4,
/* out0392_em-eta12-phi19*/	8,34,1,4,34,2,15,35,0,9,35,1,1,35,4,4,12,0,7,12,1,1,12,2,1,
/* out0393_em-eta13-phi19*/	12,32,3,1,33,3,3,34,1,9,35,1,9,44,5,1,45,5,3,6,1,1,6,2,2,11,0,1,11,2,1,12,0,3,12,1,2,
/* out0394_em-eta14-phi19*/	7,32,0,1,32,3,12,33,3,1,44,4,1,44,5,7,6,1,4,11,0,3,
/* out0395_em-eta15-phi19*/	7,32,0,13,43,2,2,44,4,3,5,1,2,5,2,1,6,1,1,11,0,2,
/* out0396_em-eta16-phi19*/	6,32,0,1,43,2,7,43,4,1,43,5,6,5,1,4,5,2,1,
/* out0397_em-eta17-phi19*/	6,42,5,1,43,0,5,43,4,6,43,5,2,5,0,5,5,1,2,
/* out0398_em-eta18-phi19*/	5,42,4,1,42,5,1,43,0,7,43,1,2,5,0,2,
/* out0399_em-eta19-phi19*/	2,42,4,3,43,1,7,
/* out0400_em-eta0-phi20*/	1,189,0,6,
/* out0401_em-eta1-phi20*/	2,188,0,3,189,0,10,
/* out0402_em-eta2-phi20*/	3,99,2,4,188,0,13,188,1,5,
/* out0403_em-eta3-phi20*/	7,98,2,5,99,1,15,99,2,8,142,0,11,142,2,3,187,0,6,188,1,11,
/* out0404_em-eta4-phi20*/	5,98,0,9,98,1,14,98,2,11,187,0,10,187,1,7,
/* out0405_em-eta5-phi20*/	8,97,0,13,97,1,2,97,2,10,98,1,1,109,1,2,109,2,1,186,0,8,187,1,9,
/* out0406_em-eta6-phi20*/	9,96,0,4,96,2,2,97,0,3,97,1,3,108,1,6,108,2,6,15,0,1,186,0,8,186,1,16,
/* out0407_em-eta7-phi20*/	8,96,0,6,107,2,10,108,1,4,14,2,1,15,0,9,15,1,1,15,2,15,66,0,6,
/* out0408_em-eta8-phi20*/	6,107,0,2,107,1,12,107,2,3,14,0,4,14,1,4,14,2,13,
/* out0409_em-eta9-phi20*/	8,106,0,3,106,2,9,107,1,2,8,1,1,13,0,1,13,2,5,14,0,4,14,1,7,
/* out0410_em-eta10-phi20*/	4,106,0,8,106,1,3,13,0,12,13,2,1,
/* out0411_em-eta11-phi20*/	11,34,3,9,35,3,5,46,5,10,47,5,7,106,0,1,106,1,1,7,1,3,7,2,5,12,0,1,13,0,3,13,1,1,
/* out0412_em-eta12-phi20*/	9,34,0,14,34,1,1,34,3,6,45,2,2,46,4,7,46,5,1,6,2,1,7,1,6,12,0,4,
/* out0413_em-eta13-phi20*/	6,34,0,2,34,1,2,45,2,8,45,4,3,45,5,12,6,2,8,
/* out0414_em-eta14-phi20*/	8,44,4,1,44,5,8,45,0,9,45,4,3,45,5,1,6,0,1,6,1,6,6,2,1,
/* out0415_em-eta15-phi20*/	6,43,2,2,44,4,11,45,0,1,45,1,5,5,2,2,6,1,4,
/* out0416_em-eta16-phi20*/	4,43,2,5,43,3,9,43,4,2,5,2,6,
/* out0417_em-eta17-phi20*/	4,42,2,5,43,4,7,5,0,6,5,2,1,
/* out0418_em-eta18-phi20*/	4,42,1,1,42,2,6,43,0,4,43,1,2,
/* out0419_em-eta19-phi20*/	2,42,1,5,43,1,5,
/* out0420_em-eta0-phi21*/	1,189,1,6,
/* out0421_em-eta1-phi21*/	2,188,3,3,189,1,10,
/* out0422_em-eta2-phi21*/	4,99,2,2,111,0,1,188,2,5,188,3,13,
/* out0423_em-eta3-phi21*/	8,99,0,16,99,1,1,99,2,2,110,2,13,111,0,3,111,1,13,187,3,6,188,2,11,
/* out0424_em-eta4-phi21*/	7,98,0,7,109,2,9,110,0,2,110,1,16,110,2,1,187,2,7,187,3,10,
/* out0425_em-eta5-phi21*/	6,108,2,1,109,0,9,109,1,14,109,2,6,186,3,8,187,2,9,
/* out0426_em-eta6-phi21*/	10,108,0,11,108,1,2,108,2,9,119,1,1,10,0,1,10,1,2,15,0,4,15,1,1,186,2,16,186,3,8,
/* out0427_em-eta7-phi21*/	11,107,0,2,107,2,3,108,0,4,108,1,4,118,1,3,118,2,3,9,2,5,10,1,5,15,0,2,15,1,14,15,2,1,
/* out0428_em-eta8-phi21*/	7,107,0,11,117,2,3,118,1,2,9,1,11,9,2,3,14,0,6,14,2,1,
/* out0429_em-eta9-phi21*/	7,106,0,1,107,0,1,117,1,6,117,2,5,8,1,2,8,2,13,14,0,2,
/* out0430_em-eta10-phi21*/	8,47,2,16,47,3,3,47,5,1,106,0,3,117,1,4,7,2,2,8,0,1,8,1,12,
/* out0431_em-eta11-phi21*/	9,46,2,2,46,5,3,47,0,9,47,3,1,47,4,14,47,5,8,7,0,3,7,1,1,7,2,9,
/* out0432_em-eta12-phi21*/	7,45,2,2,46,4,9,46,5,2,47,0,7,47,1,12,7,0,4,7,1,6,
/* out0433_em-eta13-phi21*/	7,44,2,1,44,3,1,45,2,4,45,3,14,45,4,7,6,0,4,6,2,4,
/* out0434_em-eta14-phi21*/	5,44,1,1,44,2,13,45,0,4,45,4,3,6,0,7,
/* out0435_em-eta15-phi21*/	6,44,1,7,44,2,1,45,0,2,45,1,9,0,2,2,6,0,3,
/* out0436_em-eta16-phi21*/	5,42,3,6,43,3,7,45,1,2,0,1,3,5,2,3,
/* out0437_em-eta17-phi21*/	6,42,0,1,42,2,3,42,3,9,0,1,1,5,0,2,5,2,2,
/* out0438_em-eta18-phi21*/	3,42,0,5,42,1,4,42,2,2,
/* out0439_em-eta19-phi21*/	2,42,0,1,42,1,6,
/* out0440_em-eta0-phi22*/	1,193,0,6,
/* out0441_em-eta1-phi22*/	2,192,0,3,193,0,10,
/* out0442_em-eta2-phi22*/	2,192,0,13,192,1,5,
/* out0443_em-eta3-phi22*/	8,110,0,4,110,2,2,111,0,12,111,1,3,121,1,9,121,2,12,191,0,6,192,1,11,
/* out0444_em-eta4-phi22*/	8,109,0,1,110,0,10,120,0,1,120,1,4,120,2,14,121,1,5,191,0,10,191,1,7,
/* out0445_em-eta5-phi22*/	6,109,0,6,119,0,1,119,2,12,120,1,11,190,0,8,191,1,9,
/* out0446_em-eta6-phi22*/	8,108,0,1,118,2,2,119,0,4,119,1,15,119,2,3,10,0,5,190,0,8,190,1,16,
/* out0447_em-eta7-phi22*/	9,118,0,6,118,1,3,118,2,11,4,1,2,4,2,2,9,0,3,9,2,6,10,0,10,10,1,9,
/* out0448_em-eta8-phi22*/	9,117,0,1,117,2,5,118,0,3,118,1,8,3,2,2,4,1,1,9,0,13,9,1,4,9,2,2,
/* out0449_em-eta9-phi22*/	8,117,0,9,117,1,2,117,2,3,3,1,5,3,2,2,8,0,7,8,2,3,9,1,1,
/* out0450_em-eta10-phi22*/	7,46,3,3,47,3,10,117,0,3,117,1,4,2,2,6,8,0,8,8,1,1,
/* out0451_em-eta11-phi22*/	8,46,0,8,46,1,1,46,2,11,46,3,13,47,3,2,47,4,2,2,1,7,7,0,5,
/* out0452_em-eta12-phi22*/	6,46,0,4,46,1,15,46,2,3,47,1,4,1,2,6,7,0,4,
/* out0453_em-eta13-phi22*/	4,44,3,11,45,3,2,1,1,6,1,2,3,
/* out0454_em-eta14-phi22*/	7,44,0,14,44,1,2,44,2,1,44,3,4,0,2,2,1,1,3,6,0,1,
/* out0455_em-eta15-phi22*/	3,44,0,2,44,1,6,0,2,6,
/* out0456_em-eta16-phi22*/	2,0,1,5,0,2,1,
/* out0457_em-eta17-phi22*/	3,42,0,3,42,3,1,0,1,3,
/* out0458_em-eta18-phi22*/	1,42,0,6,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	1,193,1,6,
/* out0461_em-eta1-phi23*/	2,192,3,3,193,1,10,
/* out0462_em-eta2-phi23*/	2,192,2,5,192,3,13,
/* out0463_em-eta3-phi23*/	4,121,0,14,121,2,4,191,3,6,192,2,11,
/* out0464_em-eta4-phi23*/	6,120,0,10,120,2,2,121,0,2,121,1,2,191,2,7,191,3,10,
/* out0465_em-eta5-phi23*/	6,119,0,3,119,2,1,120,0,5,120,1,1,190,3,8,191,2,9,
/* out0466_em-eta6-phi23*/	5,119,0,8,4,0,6,4,2,1,190,2,16,190,3,8,
/* out0467_em-eta7-phi23*/	4,118,0,6,4,0,8,4,1,5,4,2,13,
/* out0468_em-eta8-phi23*/	5,118,0,1,3,0,8,3,2,10,4,0,2,4,1,8,
/* out0469_em-eta9-phi23*/	4,117,0,3,3,0,7,3,1,9,3,2,2,
/* out0470_em-eta10-phi23*/	4,2,0,4,2,2,9,3,0,1,3,1,2,
/* out0471_em-eta11-phi23*/	4,46,0,3,2,0,5,2,1,7,2,2,1,
/* out0472_em-eta12-phi23*/	5,46,0,1,1,0,3,1,2,6,2,0,7,2,1,2,
/* out0473_em-eta13-phi23*/	3,1,0,6,1,1,3,1,2,1,
/* out0474_em-eta14-phi23*/	4,0,0,1,0,2,2,1,0,7,1,1,4,
/* out0475_em-eta15-phi23*/	2,0,0,4,0,2,3,
/* out0476_em-eta16-phi23*/	2,0,0,4,0,1,1,
/* out0477_em-eta17-phi23*/	2,0,0,7,0,1,3,
/* out0478_em-eta18-phi23*/	0,
/* out0479_em-eta19-phi23*/	0
};