parameter integer matrixH [0:5852] = {
/* num inputs = 144(in0-in143) */
/* num outputs = 600(out0-out599) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1750 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	0,
/* out0006_em-eta6-phi0*/	0,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	0,
/* out0010_em-eta10-phi0*/	0,
/* out0011_em-eta11-phi0*/	0,
/* out0012_em-eta12-phi0*/	0,
/* out0013_em-eta13-phi0*/	0,
/* out0014_em-eta14-phi0*/	0,
/* out0015_em-eta15-phi0*/	0,
/* out0016_em-eta16-phi0*/	0,
/* out0017_em-eta17-phi0*/	0,
/* out0018_em-eta18-phi0*/	0,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	0,
/* out0026_em-eta6-phi1*/	0,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	0,
/* out0029_em-eta9-phi1*/	0,
/* out0030_em-eta10-phi1*/	0,
/* out0031_em-eta11-phi1*/	0,
/* out0032_em-eta12-phi1*/	0,
/* out0033_em-eta13-phi1*/	0,
/* out0034_em-eta14-phi1*/	0,
/* out0035_em-eta15-phi1*/	0,
/* out0036_em-eta16-phi1*/	1,27,0,1,
/* out0037_em-eta17-phi1*/	0,
/* out0038_em-eta18-phi1*/	0,
/* out0039_em-eta19-phi1*/	4,11,1,1,11,5,2,12,1,2,12,5,4,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	0,
/* out0046_em-eta6-phi2*/	0,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	0,
/* out0049_em-eta9-phi2*/	0,
/* out0050_em-eta10-phi2*/	1,63,0,2,
/* out0051_em-eta11-phi2*/	0,
/* out0052_em-eta12-phi2*/	2,45,0,9,45,1,1,
/* out0053_em-eta13-phi2*/	2,45,0,6,45,3,4,
/* out0054_em-eta14-phi2*/	1,27,1,2,
/* out0055_em-eta15-phi2*/	2,27,0,6,27,1,7,
/* out0056_em-eta16-phi2*/	2,27,0,9,27,3,5,
/* out0057_em-eta17-phi2*/	1,27,3,8,
/* out0058_em-eta18-phi2*/	2,12,2,7,28,3,1,
/* out0059_em-eta19-phi2*/	6,11,1,3,11,5,5,12,1,5,12,2,1,12,4,1,12,5,11,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	4,103,0,3,103,1,3,115,1,2,115,2,3,
/* out0065_em-eta5-phi3*/	3,103,0,13,103,1,1,103,2,4,
/* out0066_em-eta6-phi3*/	2,91,0,13,91,1,4,
/* out0067_em-eta7-phi3*/	4,79,0,3,79,1,3,91,0,3,91,2,4,
/* out0068_em-eta8-phi3*/	3,79,0,12,79,1,1,79,2,1,
/* out0069_em-eta9-phi3*/	4,63,0,3,63,1,3,79,0,1,79,2,3,
/* out0070_em-eta10-phi3*/	3,63,0,9,63,1,1,63,2,1,
/* out0071_em-eta11-phi3*/	4,45,1,3,46,1,8,63,0,2,63,2,3,
/* out0072_em-eta12-phi3*/	5,45,0,1,45,1,12,45,2,9,46,0,4,46,1,4,
/* out0073_em-eta13-phi3*/	4,45,2,7,45,3,10,46,3,4,46,4,4,
/* out0074_em-eta14-phi3*/	4,27,1,2,28,1,9,45,3,2,46,3,8,
/* out0075_em-eta15-phi3*/	4,27,1,5,27,2,5,28,0,4,28,1,3,
/* out0076_em-eta16-phi3*/	3,27,2,11,27,3,1,28,4,3,
/* out0077_em-eta17-phi3*/	3,27,3,2,28,3,8,28,4,1,
/* out0078_em-eta18-phi3*/	3,12,2,8,12,3,4,28,3,3,
/* out0079_em-eta19-phi3*/	6,11,1,5,11,2,4,11,5,9,12,1,9,12,4,11,12,5,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	1,127,1,2,
/* out0083_em-eta3-phi4*/	4,115,1,11,127,0,16,127,1,2,127,2,2,
/* out0084_em-eta4-phi4*/	5,103,1,6,115,1,3,115,2,13,116,0,13,116,1,2,
/* out0085_em-eta5-phi4*/	6,103,1,6,103,2,12,104,0,7,104,1,1,116,0,1,116,2,1,
/* out0086_em-eta6-phi4*/	4,91,1,12,91,2,5,92,0,1,104,0,5,
/* out0087_em-eta7-phi4*/	3,79,1,5,91,2,7,92,0,7,
/* out0088_em-eta8-phi4*/	3,79,1,7,79,2,8,80,0,1,
/* out0089_em-eta9-phi4*/	3,63,1,6,79,2,4,80,0,3,
/* out0090_em-eta10-phi4*/	2,63,1,5,63,2,6,
/* out0091_em-eta11-phi4*/	4,45,4,9,46,1,1,63,2,5,64,0,4,
/* out0092_em-eta12-phi4*/	5,45,4,6,45,5,8,46,0,12,46,1,3,46,4,1,
/* out0093_em-eta13-phi4*/	4,46,2,5,46,3,3,46,4,11,46,5,7,
/* out0094_em-eta14-phi4*/	4,27,4,9,28,1,2,46,2,9,46,3,1,
/* out0095_em-eta15-phi4*/	4,27,4,3,27,5,3,28,0,9,28,1,2,
/* out0096_em-eta16-phi4*/	3,28,0,3,28,4,10,28,5,1,
/* out0097_em-eta17-phi4*/	4,28,2,6,28,3,4,28,4,2,28,5,1,
/* out0098_em-eta18-phi4*/	4,11,3,1,12,3,11,12,4,1,28,2,3,
/* out0099_em-eta19-phi4*/	5,11,0,4,11,1,7,11,2,12,11,3,4,12,4,3,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	4,127,1,3,136,0,4,136,1,2,136,2,2,
/* out0103_em-eta3-phi5*/	8,116,1,1,127,1,9,127,2,14,128,0,9,128,1,2,136,0,10,136,1,11,136,2,9,
/* out0104_em-eta4-phi5*/	5,116,0,2,116,1,13,116,2,11,117,0,3,128,0,4,
/* out0105_em-eta5-phi5*/	5,104,0,2,104,1,15,104,2,2,116,2,4,117,0,4,
/* out0106_em-eta6-phi5*/	4,92,1,7,104,0,2,104,2,13,105,0,1,
/* out0107_em-eta7-phi5*/	3,92,0,7,92,1,5,92,2,6,
/* out0108_em-eta8-phi5*/	4,80,0,3,80,1,7,92,0,1,92,2,4,
/* out0109_em-eta9-phi5*/	3,80,0,8,80,1,1,80,2,3,
/* out0110_em-eta10-phi5*/	7,63,1,1,63,2,1,64,1,9,65,0,1,65,1,12,80,0,1,80,2,2,
/* out0111_em-eta11-phi5*/	5,64,0,11,64,1,7,64,2,13,64,3,4,65,0,1,
/* out0112_em-eta12-phi5*/	8,45,4,1,45,5,8,46,5,2,48,1,2,64,0,1,64,2,1,64,3,12,65,3,4,
/* out0113_em-eta13-phi5*/	5,46,2,2,46,5,7,47,0,2,47,1,13,48,1,1,
/* out0114_em-eta14-phi5*/	5,27,4,2,47,0,13,47,1,1,47,2,1,47,3,3,
/* out0115_em-eta15-phi5*/	4,27,4,2,27,5,11,47,0,1,47,3,5,
/* out0116_em-eta16-phi5*/	3,27,5,2,28,5,12,29,1,1,
/* out0117_em-eta17-phi5*/	3,28,2,6,28,5,1,29,0,4,
/* out0118_em-eta18-phi5*/	4,11,3,7,12,3,1,28,2,1,29,0,5,
/* out0119_em-eta19-phi5*/	2,11,0,7,11,3,4,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	9,128,0,2,128,1,14,128,2,6,129,0,2,136,0,2,136,1,3,136,2,5,137,1,1,137,2,11,
/* out0124_em-eta4-phi6*/	5,117,0,3,117,1,15,128,0,1,128,2,10,129,0,5,
/* out0125_em-eta5-phi6*/	5,104,2,1,105,0,1,105,1,6,117,0,6,117,2,13,
/* out0126_em-eta6-phi6*/	4,92,1,1,105,0,13,105,1,4,105,2,4,
/* out0127_em-eta7-phi6*/	6,92,1,3,92,2,5,93,0,6,93,1,3,105,0,1,105,2,2,
/* out0128_em-eta8-phi6*/	3,80,1,6,92,2,1,93,0,8,
/* out0129_em-eta9-phi6*/	3,80,1,2,80,2,9,81,0,2,
/* out0130_em-eta10-phi6*/	6,64,4,16,64,5,6,65,0,4,65,1,4,80,2,2,81,0,2,
/* out0131_em-eta11-phi6*/	6,64,2,2,64,5,3,65,0,10,65,2,1,65,4,15,65,5,5,
/* out0132_em-eta12-phi6*/	5,47,4,5,48,1,4,65,2,8,65,3,12,65,4,1,
/* out0133_em-eta13-phi6*/	5,47,1,2,47,2,4,47,4,1,48,0,9,48,1,9,
/* out0134_em-eta14-phi6*/	4,47,2,11,47,3,2,48,0,1,48,4,6,
/* out0135_em-eta15-phi6*/	3,30,1,1,47,3,6,48,3,10,
/* out0136_em-eta16-phi6*/	3,28,5,1,29,1,8,30,1,6,
/* out0137_em-eta17-phi6*/	3,29,0,2,29,1,7,29,2,3,
/* out0138_em-eta18-phi6*/	3,29,0,5,29,2,1,29,3,5,
/* out0139_em-eta19-phi6*/	2,11,0,5,29,3,5,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	3,137,2,1,138,0,1,138,1,1,
/* out0143_em-eta3-phi7*/	7,129,0,1,129,1,14,137,1,15,137,2,4,138,0,14,138,1,1,138,2,5,
/* out0144_em-eta4-phi7*/	7,117,1,1,117,2,1,118,0,1,118,1,6,129,0,8,129,1,2,129,2,15,
/* out0145_em-eta5-phi7*/	5,105,1,2,117,2,2,118,0,15,118,1,4,118,2,4,
/* out0146_em-eta6-phi7*/	5,105,1,4,105,2,9,106,0,7,106,1,2,118,2,1,
/* out0147_em-eta7-phi7*/	4,93,1,13,93,2,2,105,2,1,106,0,3,
/* out0148_em-eta8-phi7*/	3,81,1,2,93,0,2,93,2,12,
/* out0149_em-eta9-phi7*/	3,81,0,6,81,1,7,81,2,1,
/* out0150_em-eta10-phi7*/	3,64,5,4,81,0,6,81,2,3,
/* out0151_em-eta11-phi7*/	6,64,5,3,65,2,2,65,5,11,66,0,1,66,1,13,67,1,4,
/* out0152_em-eta12-phi7*/	5,47,4,6,65,2,5,66,0,15,66,1,2,66,3,2,
/* out0153_em-eta13-phi7*/	5,47,4,4,47,5,13,48,0,6,48,5,1,66,3,1,
/* out0154_em-eta14-phi7*/	4,48,2,3,48,3,1,48,4,10,48,5,7,
/* out0155_em-eta15-phi7*/	4,29,4,4,30,1,1,48,2,8,48,3,5,
/* out0156_em-eta16-phi7*/	3,29,4,2,30,0,4,30,1,8,
/* out0157_em-eta17-phi7*/	3,29,2,7,30,0,5,30,4,1,
/* out0158_em-eta18-phi7*/	4,29,2,5,29,3,2,30,3,1,30,4,3,
/* out0159_em-eta19-phi7*/	2,29,3,4,30,3,5,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	6,130,1,7,138,0,1,138,1,14,138,2,11,139,0,2,139,2,6,
/* out0164_em-eta4-phi8*/	5,118,1,3,129,2,1,130,0,16,130,1,6,130,2,8,
/* out0165_em-eta5-phi8*/	5,106,1,1,118,1,3,118,2,11,119,0,10,119,1,3,
/* out0166_em-eta6-phi8*/	4,106,0,3,106,1,13,106,2,6,119,0,1,
/* out0167_em-eta7-phi8*/	5,93,2,1,94,0,1,94,1,6,106,0,3,106,2,7,
/* out0168_em-eta8-phi8*/	4,81,1,1,93,2,1,94,0,13,94,1,1,
/* out0169_em-eta9-phi8*/	4,81,1,6,81,2,5,82,0,1,94,0,2,
/* out0170_em-eta10-phi8*/	4,66,4,8,67,1,1,81,2,7,82,0,1,
/* out0171_em-eta11-phi8*/	7,66,1,1,66,2,5,66,4,4,66,5,1,67,0,13,67,1,11,67,4,1,
/* out0172_em-eta12-phi8*/	4,66,2,11,66,3,7,67,3,4,67,4,7,
/* out0173_em-eta13-phi8*/	6,47,5,3,48,5,3,49,1,3,50,1,4,66,3,6,67,3,6,
/* out0174_em-eta14-phi8*/	4,48,2,3,48,5,5,49,0,4,49,1,9,
/* out0175_em-eta15-phi8*/	3,29,4,5,48,2,2,49,0,10,
/* out0176_em-eta16-phi8*/	3,29,4,5,29,5,7,30,0,2,
/* out0177_em-eta17-phi8*/	4,29,5,1,30,0,5,30,4,6,30,5,1,
/* out0178_em-eta18-phi8*/	4,30,2,1,30,3,3,30,4,6,30,5,1,
/* out0179_em-eta19-phi8*/	2,30,2,2,30,3,7,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	2,139,0,5,139,1,1,
/* out0183_em-eta3-phi9*/	5,130,1,1,131,1,3,139,0,9,139,1,15,139,2,10,
/* out0184_em-eta4-phi9*/	5,119,1,3,130,1,2,130,2,8,131,0,15,131,1,5,
/* out0185_em-eta5-phi9*/	4,119,0,3,119,1,10,119,2,13,131,0,1,
/* out0186_em-eta6-phi9*/	5,106,2,2,107,0,7,107,1,8,119,0,2,119,2,3,
/* out0187_em-eta7-phi9*/	4,94,1,8,94,2,1,106,2,1,107,0,9,
/* out0188_em-eta8-phi9*/	2,94,1,1,94,2,13,
/* out0189_em-eta9-phi9*/	3,82,0,3,82,1,8,94,2,2,
/* out0190_em-eta10-phi9*/	2,66,4,2,82,0,10,
/* out0191_em-eta11-phi9*/	6,66,4,2,66,5,15,67,0,3,67,4,3,67,5,11,82,0,1,
/* out0192_em-eta12-phi9*/	5,49,4,1,67,2,15,67,3,4,67,4,5,67,5,5,
/* out0193_em-eta13-phi9*/	5,49,4,7,50,0,2,50,1,12,67,2,1,67,3,2,
/* out0194_em-eta14-phi9*/	3,49,1,4,49,2,11,50,0,6,
/* out0195_em-eta15-phi9*/	3,49,0,2,49,2,5,49,3,11,
/* out0196_em-eta16-phi9*/	3,29,5,8,30,5,1,49,3,5,
/* out0197_em-eta17-phi9*/	1,30,5,11,
/* out0198_em-eta18-phi9*/	2,30,2,9,30,5,2,
/* out0199_em-eta19-phi9*/	1,30,2,4,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	2,140,0,1,140,1,2,
/* out0203_em-eta3-phi10*/	5,131,1,3,132,1,1,140,0,15,140,1,9,140,2,15,
/* out0204_em-eta4-phi10*/	5,120,1,3,131,1,5,131,2,15,132,0,8,132,1,2,
/* out0205_em-eta5-phi10*/	4,120,0,13,120,1,10,120,2,3,131,2,1,
/* out0206_em-eta6-phi10*/	5,107,1,8,107,2,7,108,0,2,120,0,3,120,2,2,
/* out0207_em-eta7-phi10*/	4,95,0,1,95,1,8,107,2,9,108,0,1,
/* out0208_em-eta8-phi10*/	2,95,0,13,95,1,1,
/* out0209_em-eta9-phi10*/	3,82,1,8,82,2,3,95,0,2,
/* out0210_em-eta10-phi10*/	2,68,4,2,82,2,10,
/* out0211_em-eta11-phi10*/	6,68,1,11,68,2,3,68,4,2,69,0,3,69,1,15,82,2,1,
/* out0212_em-eta12-phi10*/	5,49,4,1,68,0,15,68,1,5,68,2,5,68,3,4,
/* out0213_em-eta13-phi10*/	5,49,4,7,49,5,12,50,0,2,68,0,1,68,3,2,
/* out0214_em-eta14-phi10*/	3,50,0,6,50,4,11,50,5,4,
/* out0215_em-eta15-phi10*/	3,50,2,2,50,3,11,50,4,5,
/* out0216_em-eta16-phi10*/	3,31,1,1,32,1,8,50,3,5,
/* out0217_em-eta17-phi10*/	1,31,1,11,
/* out0218_em-eta18-phi10*/	2,31,0,9,31,1,2,
/* out0219_em-eta19-phi10*/	1,31,0,4,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	1,141,1,1,
/* out0223_em-eta3-phi11*/	6,132,1,7,140,1,5,140,2,1,141,0,16,141,1,8,141,2,12,
/* out0224_em-eta4-phi11*/	5,121,1,3,132,0,8,132,1,6,132,2,16,133,0,1,
/* out0225_em-eta5-phi11*/	5,108,1,1,120,1,3,120,2,10,121,0,11,121,1,3,
/* out0226_em-eta6-phi11*/	4,108,0,6,108,1,13,108,2,3,120,2,1,
/* out0227_em-eta7-phi11*/	5,95,1,6,95,2,1,96,0,1,108,0,7,108,2,3,
/* out0228_em-eta8-phi11*/	4,83,1,1,95,1,1,95,2,13,96,0,1,
/* out0229_em-eta9-phi11*/	4,82,2,1,83,0,5,83,1,6,95,2,2,
/* out0230_em-eta10-phi11*/	4,68,4,8,68,5,1,82,2,1,83,0,7,
/* out0231_em-eta11-phi11*/	7,68,2,1,68,4,4,68,5,11,69,0,13,69,1,1,69,4,5,69,5,1,
/* out0232_em-eta12-phi11*/	4,68,2,7,68,3,4,69,3,7,69,4,11,
/* out0233_em-eta13-phi11*/	6,49,5,4,50,5,3,51,1,3,52,1,3,68,3,6,69,3,6,
/* out0234_em-eta14-phi11*/	4,50,2,4,50,5,9,51,0,3,51,1,5,
/* out0235_em-eta15-phi11*/	3,31,4,5,50,2,10,51,0,2,
/* out0236_em-eta16-phi11*/	3,31,4,5,32,0,2,32,1,7,
/* out0237_em-eta17-phi11*/	4,31,1,1,31,2,6,32,0,5,32,1,1,
/* out0238_em-eta18-phi11*/	4,31,0,1,31,1,1,31,2,6,31,3,3,
/* out0239_em-eta19-phi11*/	2,31,0,2,31,3,7,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	2,141,1,1,142,0,1,
/* out0243_em-eta3-phi12*/	6,133,1,14,133,2,1,141,1,6,141,2,4,142,0,12,142,2,7,
/* out0244_em-eta4-phi12*/	7,121,1,6,121,2,1,122,0,1,122,1,1,133,0,15,133,1,2,133,2,8,
/* out0245_em-eta5-phi12*/	5,109,1,2,121,0,4,121,1,4,121,2,15,122,0,2,
/* out0246_em-eta6-phi12*/	5,108,1,2,108,2,7,109,0,9,109,1,4,121,0,1,
/* out0247_em-eta7-phi12*/	4,96,0,2,96,1,13,108,2,3,109,0,1,
/* out0248_em-eta8-phi12*/	3,83,1,2,96,0,12,96,2,2,
/* out0249_em-eta9-phi12*/	3,83,0,1,83,1,7,83,2,6,
/* out0250_em-eta10-phi12*/	3,71,1,4,83,0,3,83,2,6,
/* out0251_em-eta11-phi12*/	6,68,5,4,69,2,1,69,5,13,70,0,2,70,1,11,71,1,3,
/* out0252_em-eta12-phi12*/	5,51,4,6,69,2,15,69,3,2,69,5,2,70,0,5,
/* out0253_em-eta13-phi12*/	5,51,1,1,51,4,4,52,0,6,52,1,13,69,3,1,
/* out0254_em-eta14-phi12*/	4,51,0,3,51,1,7,51,2,10,51,3,1,
/* out0255_em-eta15-phi12*/	4,31,4,4,31,5,1,51,0,8,51,3,5,
/* out0256_em-eta16-phi12*/	3,31,4,2,31,5,8,32,0,4,
/* out0257_em-eta17-phi12*/	3,31,2,1,32,0,5,32,4,7,
/* out0258_em-eta18-phi12*/	4,31,2,3,31,3,1,32,3,2,32,4,5,
/* out0259_em-eta19-phi12*/	2,31,3,5,32,3,4,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	9,133,2,2,134,0,6,134,1,14,134,2,2,142,0,3,142,2,9,143,0,5,143,1,3,143,2,2,
/* out0264_em-eta4-phi13*/	5,122,1,15,122,2,3,133,2,5,134,0,10,134,2,1,
/* out0265_em-eta5-phi13*/	5,109,1,6,109,2,1,110,0,1,122,0,13,122,2,6,
/* out0266_em-eta6-phi13*/	4,97,1,1,109,0,4,109,1,4,109,2,13,
/* out0267_em-eta7-phi13*/	6,96,1,3,96,2,6,97,0,5,97,1,3,109,0,2,109,2,1,
/* out0268_em-eta8-phi13*/	3,84,1,6,96,2,8,97,0,1,
/* out0269_em-eta9-phi13*/	3,83,2,2,84,0,9,84,1,2,
/* out0270_em-eta10-phi13*/	6,70,4,16,70,5,4,71,0,4,71,1,6,83,2,2,84,0,2,
/* out0271_em-eta11-phi13*/	6,70,0,1,70,1,5,70,2,15,71,0,10,71,1,3,71,4,2,
/* out0272_em-eta12-phi13*/	5,51,4,5,51,5,4,70,0,8,70,2,1,70,3,12,
/* out0273_em-eta13-phi13*/	5,51,4,1,51,5,9,52,0,9,52,4,4,52,5,2,
/* out0274_em-eta14-phi13*/	4,51,2,6,52,0,1,52,3,2,52,4,11,
/* out0275_em-eta15-phi13*/	3,31,5,1,51,3,10,52,3,6,
/* out0276_em-eta16-phi13*/	3,31,5,6,32,5,8,33,1,1,
/* out0277_em-eta17-phi13*/	3,32,2,2,32,4,3,32,5,7,
/* out0278_em-eta18-phi13*/	3,32,2,5,32,3,5,32,4,1,
/* out0279_em-eta19-phi13*/	2,13,4,5,32,3,5,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	4,135,1,3,143,0,2,143,1,2,143,2,4,
/* out0283_em-eta3-phi14*/	8,123,1,1,134,1,2,134,2,9,135,0,14,135,1,9,143,0,9,143,1,11,143,2,10,
/* out0284_em-eta4-phi14*/	5,122,2,3,123,0,11,123,1,13,123,2,2,134,2,4,
/* out0285_em-eta5-phi14*/	5,110,0,2,110,1,15,110,2,2,122,2,4,123,0,4,
/* out0286_em-eta6-phi14*/	4,97,1,7,109,2,1,110,0,13,110,2,2,
/* out0287_em-eta7-phi14*/	3,97,0,6,97,1,5,97,2,7,
/* out0288_em-eta8-phi14*/	4,84,1,7,84,2,3,97,0,4,97,2,1,
/* out0289_em-eta9-phi14*/	3,84,0,3,84,1,1,84,2,8,
/* out0290_em-eta10-phi14*/	7,70,5,12,71,0,1,71,5,9,72,0,1,72,1,1,84,0,2,84,2,1,
/* out0291_em-eta11-phi14*/	5,71,0,1,71,2,11,71,3,4,71,4,13,71,5,7,
/* out0292_em-eta12-phi14*/	8,51,5,2,53,1,2,53,4,1,54,1,8,70,3,4,71,2,1,71,3,12,71,4,1,
/* out0293_em-eta13-phi14*/	5,51,5,1,52,2,2,52,5,13,53,0,2,53,1,7,
/* out0294_em-eta14-phi14*/	5,33,4,2,52,2,13,52,3,3,52,4,1,52,5,1,
/* out0295_em-eta15-phi14*/	4,33,4,2,34,1,11,52,2,1,52,3,5,
/* out0296_em-eta16-phi14*/	3,32,5,1,33,1,12,34,1,2,
/* out0297_em-eta17-phi14*/	3,32,2,4,33,0,6,33,1,1,
/* out0298_em-eta18-phi14*/	4,13,5,7,14,5,1,32,2,5,33,0,1,
/* out0299_em-eta19-phi14*/	2,13,4,7,13,5,4,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	1,135,1,2,
/* out0303_em-eta3-phi15*/	3,135,0,2,135,1,2,135,2,16,
/* out0304_em-eta4-phi15*/	4,111,1,6,123,1,2,123,2,13,124,2,5,
/* out0305_em-eta5-phi15*/	6,110,1,1,110,2,7,111,0,12,111,1,6,123,0,1,123,2,1,
/* out0306_em-eta6-phi15*/	4,97,2,1,98,0,5,98,1,12,110,2,5,
/* out0307_em-eta7-phi15*/	3,85,1,5,97,2,7,98,0,7,
/* out0308_em-eta8-phi15*/	3,84,2,1,85,0,8,85,1,7,
/* out0309_em-eta9-phi15*/	3,72,1,6,84,2,3,85,0,4,
/* out0310_em-eta10-phi15*/	2,72,0,6,72,1,5,
/* out0311_em-eta11-phi15*/	4,53,4,9,53,5,1,71,2,4,72,0,5,
/* out0312_em-eta12-phi15*/	5,53,2,1,53,4,6,53,5,3,54,0,12,54,1,8,
/* out0313_em-eta13-phi15*/	4,53,0,5,53,1,7,53,2,11,53,3,3,
/* out0314_em-eta14-phi15*/	4,33,4,9,33,5,2,53,0,9,53,3,1,
/* out0315_em-eta15-phi15*/	4,33,4,3,33,5,2,34,0,9,34,1,3,
/* out0316_em-eta16-phi15*/	3,33,1,1,33,2,10,34,0,3,
/* out0317_em-eta17-phi15*/	4,33,0,6,33,1,1,33,2,2,33,3,4,
/* out0318_em-eta18-phi15*/	4,13,5,1,14,4,1,14,5,11,33,0,3,
/* out0319_em-eta19-phi15*/	5,13,4,4,13,5,4,14,0,12,14,1,7,14,4,3,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	1,125,1,2,
/* out0323_em-eta3-phi16*/	4,124,1,8,124,2,3,125,0,10,125,1,10,
/* out0324_em-eta4-phi16*/	6,111,1,3,111,2,3,112,0,6,112,1,9,124,1,8,124,2,8,
/* out0325_em-eta5-phi16*/	5,99,1,7,111,0,4,111,1,1,111,2,13,112,0,2,
/* out0326_em-eta6-phi16*/	4,86,1,1,98,1,4,98,2,13,99,0,5,
/* out0327_em-eta7-phi16*/	6,85,1,3,85,2,3,86,0,3,86,1,3,98,0,4,98,2,3,
/* out0328_em-eta8-phi16*/	5,73,1,1,85,0,1,85,1,1,85,2,12,86,0,1,
/* out0329_em-eta9-phi16*/	6,72,1,3,72,2,3,73,0,2,73,1,1,85,0,3,85,2,1,
/* out0330_em-eta10-phi16*/	3,72,0,1,72,1,1,72,2,9,
/* out0331_em-eta11-phi16*/	6,53,5,8,54,5,3,55,1,2,56,1,3,72,0,3,72,2,2,
/* out0332_em-eta12-phi16*/	5,53,5,4,54,0,4,54,2,1,54,4,9,54,5,12,
/* out0333_em-eta13-phi16*/	4,53,2,4,53,3,4,54,3,10,54,4,7,
/* out0334_em-eta14-phi16*/	4,33,5,9,34,5,2,53,3,8,54,3,2,
/* out0335_em-eta15-phi16*/	4,33,5,3,34,0,4,34,4,5,34,5,5,
/* out0336_em-eta16-phi16*/	3,33,2,3,34,3,1,34,4,11,
/* out0337_em-eta17-phi16*/	3,33,2,1,33,3,8,34,3,2,
/* out0338_em-eta18-phi16*/	3,14,2,8,14,5,4,33,3,3,
/* out0339_em-eta19-phi16*/	6,13,1,9,13,3,9,14,0,4,14,1,5,14,3,1,14,4,11,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	5,125,1,2,125,2,1,126,0,4,126,1,2,126,2,2,
/* out0343_em-eta3-phi17*/	9,112,1,1,113,0,2,113,1,9,125,0,6,125,1,2,125,2,15,126,0,10,126,1,11,126,2,9,
/* out0344_em-eta4-phi17*/	5,100,1,3,112,0,4,112,1,6,112,2,15,113,0,5,
/* out0345_em-eta5-phi17*/	7,99,0,1,99,1,9,99,2,10,100,0,2,100,1,1,112,0,4,112,2,1,
/* out0346_em-eta6-phi17*/	5,86,1,6,86,2,2,87,1,1,99,0,10,99,2,5,
/* out0347_em-eta7-phi17*/	3,86,0,7,86,1,6,86,2,6,
/* out0348_em-eta8-phi17*/	2,73,1,10,86,0,5,
/* out0349_em-eta9-phi17*/	3,73,0,8,73,1,3,73,2,1,
/* out0350_em-eta10-phi17*/	6,55,4,16,55,5,4,56,0,1,56,1,1,72,2,2,73,0,3,
/* out0351_em-eta11-phi17*/	4,55,1,9,55,2,6,56,0,8,56,1,12,
/* out0352_em-eta12-phi17*/	6,35,4,2,54,2,9,54,5,1,55,0,12,55,1,5,55,2,1,
/* out0353_em-eta13-phi17*/	4,35,4,8,36,1,8,54,2,6,54,3,4,
/* out0354_em-eta14-phi17*/	3,34,5,2,35,1,11,36,1,7,
/* out0355_em-eta15-phi17*/	4,34,2,6,34,5,7,35,0,3,35,1,2,
/* out0356_em-eta16-phi17*/	2,34,2,9,34,3,5,
/* out0357_em-eta17-phi17*/	2,16,1,4,34,3,8,
/* out0358_em-eta18-phi17*/	4,14,2,7,15,1,3,16,1,1,33,3,1,
/* out0359_em-eta19-phi17*/	6,13,1,5,13,3,5,14,1,3,14,2,1,14,3,11,14,4,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	9,101,1,2,113,0,2,113,1,7,113,2,13,114,0,11,114,2,1,126,0,2,126,1,3,126,2,5,
/* out0364_em-eta4-phi18*/	6,100,1,11,100,2,7,101,0,2,101,1,3,113,0,7,113,2,3,
/* out0365_em-eta5-phi18*/	6,87,1,6,87,2,1,99,2,1,100,0,14,100,1,1,100,2,5,
/* out0366_em-eta6-phi18*/	4,86,2,1,87,0,10,87,1,9,87,2,2,
/* out0367_em-eta7-phi18*/	3,74,1,9,86,2,7,87,0,3,
/* out0368_em-eta8-phi18*/	4,73,1,1,73,2,6,74,0,7,74,1,2,
/* out0369_em-eta9-phi18*/	3,57,1,2,73,0,1,73,2,9,
/* out0370_em-eta10-phi18*/	7,55,5,12,56,0,3,56,4,1,56,5,14,57,0,1,57,1,1,73,0,2,
/* out0371_em-eta11-phi18*/	6,55,2,8,56,0,4,56,2,1,56,3,5,56,4,15,56,5,2,
/* out0372_em-eta12-phi18*/	6,35,4,3,35,5,6,55,0,4,55,2,1,55,3,15,56,3,2,
/* out0373_em-eta13-phi18*/	5,35,4,3,35,5,8,36,0,12,36,1,1,36,4,2,
/* out0374_em-eta14-phi18*/	4,35,1,2,35,2,13,36,0,4,36,4,1,
/* out0375_em-eta15-phi18*/	4,15,4,1,35,0,13,35,1,1,35,3,3,
/* out0376_em-eta16-phi18*/	3,15,4,13,16,1,1,34,2,1,
/* out0377_em-eta17-phi18*/	2,16,0,3,16,1,9,
/* out0378_em-eta18-phi18*/	3,15,1,9,15,2,1,16,1,1,
/* out0379_em-eta19-phi18*/	6,13,1,2,13,3,2,14,1,1,14,3,4,15,0,4,15,1,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	3,102,0,1,102,1,1,114,0,1,
/* out0383_em-eta3-phi19*/	7,101,1,8,101,2,7,102,0,14,102,1,1,102,2,5,114,0,4,114,2,15,
/* out0384_em-eta4-phi19*/	6,88,1,6,88,2,1,100,2,2,101,0,14,101,1,3,101,2,8,
/* out0385_em-eta5-phi19*/	5,87,2,2,88,0,11,88,1,10,88,2,2,100,2,2,
/* out0386_em-eta6-phi19*/	5,75,0,1,75,1,8,87,0,2,87,2,11,88,0,2,
/* out0387_em-eta7-phi19*/	4,74,1,5,74,2,9,75,0,3,87,0,1,
/* out0388_em-eta8-phi19*/	3,57,1,2,74,0,9,74,2,4,
/* out0389_em-eta9-phi19*/	3,57,0,1,57,1,11,57,2,1,
/* out0390_em-eta10-phi19*/	2,56,2,4,57,0,10,
/* out0391_em-eta11-phi19*/	4,37,4,12,38,1,6,56,2,11,56,3,5,
/* out0392_em-eta12-phi19*/	6,35,5,2,36,5,4,37,1,10,38,1,9,55,3,1,56,3,4,
/* out0393_em-eta13-phi19*/	4,36,2,6,36,4,6,36,5,12,37,0,1,
/* out0394_em-eta14-phi19*/	4,35,2,3,35,3,2,36,3,9,36,4,7,
/* out0395_em-eta15-phi19*/	4,15,4,1,15,5,5,35,3,11,36,3,1,
/* out0396_em-eta16-phi19*/	3,15,4,1,15,5,9,16,0,4,
/* out0397_em-eta17-phi19*/	3,15,2,3,16,0,9,16,4,1,
/* out0398_em-eta18-phi19*/	3,15,0,1,15,1,2,15,2,8,
/* out0399_em-eta19-phi19*/	2,15,0,8,15,3,1,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	7,89,1,5,89,2,2,90,0,2,90,2,6,102,0,1,102,1,14,102,2,11,
/* out0404_em-eta4-phi20*/	5,88,2,2,89,0,14,89,1,11,89,2,5,101,2,1,
/* out0405_em-eta5-phi20*/	5,75,1,1,76,0,3,76,1,9,88,0,3,88,2,11,
/* out0406_em-eta6-phi20*/	4,75,0,2,75,1,7,75,2,12,76,0,1,
/* out0407_em-eta7-phi20*/	3,58,1,7,74,2,2,75,0,10,
/* out0408_em-eta8-phi20*/	4,57,2,1,58,0,6,58,1,7,74,2,1,
/* out0409_em-eta9-phi20*/	3,39,1,1,57,2,11,58,0,2,
/* out0410_em-eta10-phi20*/	6,37,4,1,37,5,6,38,5,3,39,1,1,57,0,4,57,2,3,
/* out0411_em-eta11-phi20*/	6,37,4,3,37,5,10,38,0,13,38,1,1,38,4,6,38,5,3,
/* out0412_em-eta12-phi20*/	6,37,0,3,37,1,6,37,2,14,37,3,3,38,0,3,38,4,1,
/* out0413_em-eta13-phi20*/	3,17,4,7,36,2,7,37,0,11,
/* out0414_em-eta14-phi20*/	4,17,4,4,18,1,9,36,2,3,36,3,4,
/* out0415_em-eta15-phi20*/	5,15,5,1,16,5,4,17,1,6,18,1,4,36,3,2,
/* out0416_em-eta16-phi20*/	3,15,5,1,16,4,2,16,5,12,
/* out0417_em-eta17-phi20*/	2,16,3,1,16,4,11,
/* out0418_em-eta18-phi20*/	4,15,2,4,15,3,4,16,3,1,16,4,2,
/* out0419_em-eta19-phi20*/	2,15,0,3,15,3,6,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	2,90,0,5,90,1,1,
/* out0423_em-eta3-phi21*/	5,77,1,3,89,2,1,90,0,9,90,1,15,90,2,10,
/* out0424_em-eta4-phi21*/	6,76,1,2,76,2,1,77,0,7,77,1,13,89,0,2,89,2,8,
/* out0425_em-eta5-phi21*/	4,76,0,7,76,1,5,76,2,15,77,0,1,
/* out0426_em-eta6-phi21*/	3,59,1,14,75,2,3,76,0,5,
/* out0427_em-eta7-phi21*/	5,58,1,2,58,2,7,59,0,8,59,1,2,75,2,1,
/* out0428_em-eta8-phi21*/	2,58,0,6,58,2,9,
/* out0429_em-eta9-phi21*/	2,39,1,11,58,0,2,
/* out0430_em-eta10-phi21*/	3,38,5,2,39,0,7,39,1,3,
/* out0431_em-eta11-phi21*/	5,38,2,16,38,3,3,38,4,5,38,5,8,39,0,1,
/* out0432_em-eta12-phi21*/	5,17,5,1,37,2,2,37,3,11,38,3,13,38,4,4,
/* out0433_em-eta13-phi21*/	5,17,4,4,17,5,15,18,0,2,37,0,1,37,3,2,
/* out0434_em-eta14-phi21*/	4,17,2,3,17,4,1,18,0,14,18,1,3,
/* out0435_em-eta15-phi21*/	3,17,0,3,17,1,10,17,2,5,
/* out0436_em-eta16-phi21*/	2,16,2,9,17,0,5,
/* out0437_em-eta17-phi21*/	2,16,2,7,16,3,5,
/* out0438_em-eta18-phi21*/	2,15,3,1,16,3,9,
/* out0439_em-eta19-phi21*/	1,15,3,4,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	1,78,1,2,
/* out0443_em-eta3-phi22*/	5,61,1,1,77,2,3,78,0,16,78,1,13,78,2,10,
/* out0444_em-eta4-phi22*/	6,60,1,1,60,2,2,61,0,2,61,1,8,77,0,7,77,2,13,
/* out0445_em-eta5-phi22*/	4,60,0,7,60,1,15,60,2,5,77,0,1,
/* out0446_em-eta6-phi22*/	3,41,1,3,59,2,14,60,0,5,
/* out0447_em-eta7-phi22*/	5,40,1,7,40,2,2,41,1,1,59,0,8,59,2,2,
/* out0448_em-eta8-phi22*/	2,40,0,6,40,1,9,
/* out0449_em-eta9-phi22*/	2,39,2,11,40,0,2,
/* out0450_em-eta10-phi22*/	3,19,5,2,39,0,7,39,2,3,
/* out0451_em-eta11-phi22*/	5,19,4,16,19,5,8,20,0,5,20,1,3,39,0,1,
/* out0452_em-eta12-phi22*/	5,18,5,1,19,1,11,19,2,2,20,0,4,20,1,13,
/* out0453_em-eta13-phi22*/	5,18,2,4,18,4,2,18,5,15,19,0,1,19,1,2,
/* out0454_em-eta14-phi22*/	4,17,2,3,18,2,1,18,3,3,18,4,14,
/* out0455_em-eta15-phi22*/	3,17,0,3,17,2,5,17,3,10,
/* out0456_em-eta16-phi22*/	2,0,4,9,17,0,5,
/* out0457_em-eta17-phi22*/	2,0,4,7,1,1,5,
/* out0458_em-eta18-phi22*/	2,0,1,1,1,1,9,
/* out0459_em-eta19-phi22*/	1,0,1,4,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	1,62,1,1,
/* out0463_em-eta3-phi23*/	7,61,1,2,61,2,5,62,0,16,62,1,8,62,2,12,78,1,1,78,2,6,
/* out0464_em-eta4-phi23*/	5,42,1,2,43,1,1,61,0,14,61,1,5,61,2,11,
/* out0465_em-eta5-phi23*/	5,41,2,1,42,0,3,42,1,11,60,0,3,60,2,9,
/* out0466_em-eta6-phi23*/	4,41,0,2,41,1,12,41,2,7,60,0,1,
/* out0467_em-eta7-phi23*/	3,22,1,2,40,2,7,41,0,10,
/* out0468_em-eta8-phi23*/	4,21,1,1,22,1,1,40,0,6,40,2,7,
/* out0469_em-eta9-phi23*/	3,21,1,11,39,2,1,40,0,2,
/* out0470_em-eta10-phi23*/	6,19,5,3,20,2,1,20,5,6,21,0,4,21,1,3,39,2,1,
/* out0471_em-eta11-phi23*/	6,19,5,3,20,0,6,20,2,3,20,3,1,20,4,13,20,5,10,
/* out0472_em-eta12-phi23*/	6,19,0,3,19,1,3,19,2,14,19,3,6,20,0,1,20,4,3,
/* out0473_em-eta13-phi23*/	3,2,4,7,18,2,7,19,0,11,
/* out0474_em-eta14-phi23*/	4,2,4,3,3,1,4,18,2,4,18,3,9,
/* out0475_em-eta15-phi23*/	5,0,5,4,1,5,1,3,1,2,17,3,6,18,3,4,
/* out0476_em-eta16-phi23*/	3,0,5,12,1,0,2,1,5,1,
/* out0477_em-eta17-phi23*/	2,1,0,11,1,1,1,
/* out0478_em-eta18-phi23*/	4,0,1,4,0,2,4,1,0,2,1,1,1,
/* out0479_em-eta19-phi23*/	2,0,0,3,0,1,6,
/* out0480_em-eta0-phi24*/	0,
/* out0481_em-eta1-phi24*/	0,
/* out0482_em-eta2-phi24*/	2,44,0,1,62,1,1,
/* out0483_em-eta3-phi24*/	6,43,1,7,43,2,8,44,0,12,44,2,7,62,1,6,62,2,4,
/* out0484_em-eta4-phi24*/	6,24,1,2,42,1,1,42,2,6,43,0,14,43,1,8,43,2,3,
/* out0485_em-eta5-phi24*/	5,23,1,2,24,1,2,42,0,11,42,1,2,42,2,10,
/* out0486_em-eta6-phi24*/	5,23,0,2,23,1,11,41,0,1,41,2,8,42,0,2,
/* out0487_em-eta7-phi24*/	4,22,1,9,22,2,5,23,0,1,41,0,3,
/* out0488_em-eta8-phi24*/	3,21,2,2,22,0,9,22,1,4,
/* out0489_em-eta9-phi24*/	3,21,0,1,21,1,1,21,2,11,
/* out0490_em-eta10-phi24*/	2,4,4,4,21,0,10,
/* out0491_em-eta11-phi24*/	4,4,4,11,5,1,5,20,2,12,20,3,6,
/* out0492_em-eta12-phi24*/	6,2,5,4,3,5,2,4,1,1,5,1,4,19,3,10,20,3,9,
/* out0493_em-eta13-phi24*/	4,2,4,6,2,5,12,3,0,6,19,0,1,
/* out0494_em-eta14-phi24*/	4,2,1,2,2,2,3,3,0,7,3,1,9,
/* out0495_em-eta15-phi24*/	4,1,2,1,1,5,5,2,1,11,3,1,1,
/* out0496_em-eta16-phi24*/	3,1,2,1,1,4,4,1,5,9,
/* out0497_em-eta17-phi24*/	3,0,2,3,1,0,1,1,4,9,
/* out0498_em-eta18-phi24*/	3,0,0,1,0,2,8,0,3,2,
/* out0499_em-eta19-phi24*/	2,0,0,8,0,1,1,
/* out0500_em-eta0-phi25*/	0,
/* out0501_em-eta1-phi25*/	0,
/* out0502_em-eta2-phi25*/	0,
/* out0503_em-eta3-phi25*/	9,25,0,2,25,1,13,25,2,7,26,0,5,26,1,3,26,2,2,43,2,2,44,0,3,44,2,9,
/* out0504_em-eta4-phi25*/	6,24,1,7,24,2,11,25,0,7,25,1,3,43,0,2,43,2,3,
/* out0505_em-eta5-phi25*/	6,8,1,1,23,1,1,23,2,6,24,0,14,24,1,5,24,2,1,
/* out0506_em-eta6-phi25*/	4,7,1,1,23,0,10,23,1,2,23,2,9,
/* out0507_em-eta7-phi25*/	3,7,1,7,22,2,9,23,0,3,
/* out0508_em-eta8-phi25*/	4,6,1,6,6,2,1,22,0,7,22,2,2,
/* out0509_em-eta9-phi25*/	3,6,0,1,6,1,9,21,2,2,
/* out0510_em-eta10-phi25*/	7,4,5,14,5,0,1,5,4,3,5,5,12,6,0,2,21,0,1,21,2,1,
/* out0511_em-eta11-phi25*/	6,4,2,8,4,4,1,4,5,2,5,0,15,5,1,5,5,4,4,
/* out0512_em-eta12-phi25*/	6,3,2,3,3,5,6,4,0,4,4,1,15,4,2,1,5,1,2,
/* out0513_em-eta13-phi25*/	5,3,0,2,3,2,3,3,3,1,3,4,12,3,5,8,
/* out0514_em-eta14-phi25*/	4,2,2,13,2,3,2,3,0,1,3,4,4,
/* out0515_em-eta15-phi25*/	4,1,2,1,2,0,13,2,1,3,2,3,1,
/* out0516_em-eta16-phi25*/	2,1,2,13,1,3,1,
/* out0517_em-eta17-phi25*/	2,1,3,9,1,4,3,
/* out0518_em-eta18-phi25*/	3,0,2,1,0,3,9,1,3,1,
/* out0519_em-eta19-phi25*/	2,0,0,4,0,3,2,
/* out0520_em-eta0-phi26*/	0,
/* out0521_em-eta1-phi26*/	0,
/* out0522_em-eta2-phi26*/	5,10,1,1,10,2,2,26,0,2,26,1,2,26,2,4,
/* out0523_em-eta3-phi26*/	9,9,2,1,10,0,6,10,1,15,10,2,2,25,0,2,25,2,9,26,0,9,26,1,11,26,2,10,
/* out0524_em-eta4-phi26*/	5,9,0,4,9,1,15,9,2,6,24,2,3,25,0,5,
/* out0525_em-eta5-phi26*/	7,8,0,1,8,1,10,8,2,9,9,0,4,9,1,1,24,0,2,24,2,1,
/* out0526_em-eta6-phi26*/	5,7,1,2,7,2,6,8,0,10,8,1,5,23,2,1,
/* out0527_em-eta7-phi26*/	3,7,0,7,7,1,6,7,2,6,
/* out0528_em-eta8-phi26*/	2,6,2,10,7,0,5,
/* out0529_em-eta9-phi26*/	3,6,0,8,6,1,1,6,2,3,
/* out0530_em-eta10-phi26*/	5,5,2,16,5,3,1,5,4,1,5,5,4,6,0,3,
/* out0531_em-eta11-phi26*/	4,4,2,6,4,3,9,5,3,12,5,4,8,
/* out0532_em-eta12-phi26*/	4,3,2,2,4,0,12,4,2,1,4,3,5,
/* out0533_em-eta13-phi26*/	2,3,2,8,3,3,8,
/* out0534_em-eta14-phi26*/	2,2,3,11,3,3,7,
/* out0535_em-eta15-phi26*/	2,2,0,3,2,3,2,
/* out0536_em-eta16-phi26*/	0,
/* out0537_em-eta17-phi26*/	1,1,3,4,
/* out0538_em-eta18-phi26*/	2,0,3,3,1,3,1,
/* out0539_em-eta19-phi26*/	0,
/* out0540_em-eta0-phi27*/	0,
/* out0541_em-eta1-phi27*/	0,
/* out0542_em-eta2-phi27*/	1,10,2,2,
/* out0543_em-eta3-phi27*/	2,10,0,10,10,2,10,
/* out0544_em-eta4-phi27*/	2,9,0,6,9,2,9,
/* out0545_em-eta5-phi27*/	2,8,2,7,9,0,2,
/* out0546_em-eta6-phi27*/	2,7,2,1,8,0,5,
/* out0547_em-eta7-phi27*/	2,7,0,3,7,2,3,
/* out0548_em-eta8-phi27*/	2,6,2,1,7,0,1,
/* out0549_em-eta9-phi27*/	2,6,0,2,6,2,1,
/* out0550_em-eta10-phi27*/	0,
/* out0551_em-eta11-phi27*/	2,4,3,2,5,3,3,
/* out0552_em-eta12-phi27*/	0,
/* out0553_em-eta13-phi27*/	0,
/* out0554_em-eta14-phi27*/	0,
/* out0555_em-eta15-phi27*/	0,
/* out0556_em-eta16-phi27*/	0,
/* out0557_em-eta17-phi27*/	0,
/* out0558_em-eta18-phi27*/	0,
/* out0559_em-eta19-phi27*/	0,
/* out0560_em-eta0-phi28*/	0,
/* out0561_em-eta1-phi28*/	0,
/* out0562_em-eta2-phi28*/	0,
/* out0563_em-eta3-phi28*/	0,
/* out0564_em-eta4-phi28*/	0,
/* out0565_em-eta5-phi28*/	0,
/* out0566_em-eta6-phi28*/	0,
/* out0567_em-eta7-phi28*/	0,
/* out0568_em-eta8-phi28*/	0,
/* out0569_em-eta9-phi28*/	0,
/* out0570_em-eta10-phi28*/	0,
/* out0571_em-eta11-phi28*/	0,
/* out0572_em-eta12-phi28*/	0,
/* out0573_em-eta13-phi28*/	0,
/* out0574_em-eta14-phi28*/	0,
/* out0575_em-eta15-phi28*/	0,
/* out0576_em-eta16-phi28*/	0,
/* out0577_em-eta17-phi28*/	0,
/* out0578_em-eta18-phi28*/	0,
/* out0579_em-eta19-phi28*/	0,
/* out0580_em-eta0-phi29*/	0,
/* out0581_em-eta1-phi29*/	0,
/* out0582_em-eta2-phi29*/	0,
/* out0583_em-eta3-phi29*/	0,
/* out0584_em-eta4-phi29*/	0,
/* out0585_em-eta5-phi29*/	0,
/* out0586_em-eta6-phi29*/	0,
/* out0587_em-eta7-phi29*/	0,
/* out0588_em-eta8-phi29*/	0,
/* out0589_em-eta9-phi29*/	0,
/* out0590_em-eta10-phi29*/	0,
/* out0591_em-eta11-phi29*/	0,
/* out0592_em-eta12-phi29*/	0,
/* out0593_em-eta13-phi29*/	0,
/* out0594_em-eta14-phi29*/	0,
/* out0595_em-eta15-phi29*/	0,
/* out0596_em-eta16-phi29*/	0,
/* out0597_em-eta17-phi29*/	0,
/* out0598_em-eta18-phi29*/	0,
/* out0599_em-eta19-phi29*/	0
};