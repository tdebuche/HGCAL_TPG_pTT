parameter integer matrixH [0:5183] = {
/* num inputs = 100(in0-in99) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 10 */
//* total number of input in adders 1567 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	4,75,0,2,75,1,6,85,1,9,85,2,15,
/* out0006_em-eta6-phi0*/	3,75,0,14,75,1,2,75,2,7,
/* out0007_em-eta7-phi0*/	3,65,0,12,65,1,6,65,2,1,
/* out0008_em-eta8-phi0*/	4,54,0,2,54,1,3,65,0,4,65,2,4,
/* out0009_em-eta9-phi0*/	2,54,0,12,54,1,1,
/* out0010_em-eta10-phi0*/	4,43,0,2,43,1,1,54,0,2,54,2,2,
/* out0011_em-eta11-phi0*/	2,43,0,9,104,0,9,
/* out0012_em-eta12-phi0*/	6,32,1,1,43,0,3,43,2,1,104,0,6,104,1,3,104,2,7,
/* out0013_em-eta13-phi0*/	3,32,0,5,96,0,4,104,2,8,
/* out0014_em-eta14-phi0*/	4,32,0,5,96,0,10,96,1,1,96,2,2,
/* out0015_em-eta15-phi0*/	2,32,0,1,96,2,8,
/* out0016_em-eta16-phi0*/	3,22,0,3,88,0,8,96,2,3,
/* out0017_em-eta17-phi0*/	3,22,0,3,88,0,4,88,2,2,
/* out0018_em-eta18-phi0*/	2,22,0,1,88,2,5,
/* out0019_em-eta19-phi0*/	1,88,2,2,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	1,86,1,2,
/* out0025_em-eta5-phi1*/	6,75,1,4,85,1,7,85,2,1,86,0,15,86,1,5,86,2,3,
/* out0026_em-eta6-phi1*/	6,75,1,4,75,2,9,76,0,9,76,1,2,86,0,1,86,2,2,
/* out0027_em-eta7-phi1*/	4,65,1,10,65,2,5,66,0,1,76,0,5,
/* out0028_em-eta8-phi1*/	3,54,1,6,65,2,6,66,0,6,
/* out0029_em-eta9-phi1*/	2,54,1,6,54,2,9,
/* out0030_em-eta10-phi1*/	3,43,1,8,54,2,4,55,0,1,
/* out0031_em-eta11-phi1*/	6,43,0,2,43,1,4,43,2,5,104,0,1,104,1,2,111,2,8,
/* out0032_em-eta12-phi1*/	6,32,1,3,43,2,6,104,1,9,105,0,3,111,1,1,111,2,2,
/* out0033_em-eta13-phi1*/	8,32,0,2,32,1,5,96,0,1,96,1,1,104,1,2,104,2,1,105,0,3,105,2,3,
/* out0034_em-eta14-phi1*/	5,32,0,3,32,2,4,96,0,1,96,1,8,105,2,1,
/* out0035_em-eta15-phi1*/	5,22,1,3,32,2,2,96,1,5,96,2,2,97,0,1,
/* out0036_em-eta16-phi1*/	5,22,0,3,22,1,1,88,0,3,88,1,3,96,2,1,
/* out0037_em-eta17-phi1*/	4,22,0,4,88,0,1,88,1,5,88,2,1,
/* out0038_em-eta18-phi1*/	4,22,0,2,22,2,1,88,1,2,88,2,3,
/* out0039_em-eta19-phi1*/	2,22,2,1,88,2,2,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	4,86,1,1,94,0,4,94,1,1,94,2,2,
/* out0045_em-eta5-phi2*/	7,86,1,8,86,2,10,87,0,7,87,1,2,94,0,11,94,1,12,94,2,10,
/* out0046_em-eta6-phi2*/	5,76,0,1,76,1,14,76,2,6,86,2,1,87,0,6,
/* out0047_em-eta7-phi2*/	5,66,0,1,66,1,10,76,0,1,76,2,10,77,0,2,
/* out0048_em-eta8-phi2*/	3,66,0,7,66,1,4,66,2,8,
/* out0049_em-eta9-phi2*/	5,54,2,1,55,0,5,55,1,7,66,0,1,66,2,3,
/* out0050_em-eta10-phi2*/	3,43,1,1,55,0,10,55,2,2,
/* out0051_em-eta11-phi2*/	7,43,1,2,43,2,3,44,0,3,44,1,1,55,2,1,111,1,8,111,2,6,
/* out0052_em-eta12-phi2*/	6,32,1,2,43,2,1,44,0,6,105,0,7,105,1,2,111,1,5,
/* out0053_em-eta13-phi2*/	6,32,1,5,32,2,2,44,0,1,105,0,3,105,1,2,105,2,5,
/* out0054_em-eta14-phi2*/	4,32,2,6,96,1,1,97,0,3,105,2,5,
/* out0055_em-eta15-phi2*/	4,22,1,4,32,2,1,97,0,7,97,2,1,
/* out0056_em-eta16-phi2*/	3,22,1,4,88,1,1,97,2,6,
/* out0057_em-eta17-phi2*/	4,22,2,3,88,1,3,89,1,1,97,2,1,
/* out0058_em-eta18-phi2*/	3,22,2,3,88,1,2,89,1,2,
/* out0059_em-eta19-phi2*/	2,88,2,1,89,1,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	2,95,0,4,95,1,2,
/* out0065_em-eta5-phi3*/	10,87,0,1,87,1,14,87,2,5,88,0,1,94,0,1,94,1,3,94,2,4,95,0,12,95,1,2,95,2,8,
/* out0066_em-eta6-phi3*/	5,77,0,2,77,1,11,87,0,2,87,2,11,88,0,2,
/* out0067_em-eta7-phi3*/	4,66,1,1,77,0,12,77,1,2,77,2,8,
/* out0068_em-eta8-phi3*/	4,66,1,1,66,2,5,67,0,9,67,1,3,
/* out0069_em-eta9-phi3*/	3,55,1,9,55,2,1,67,0,5,
/* out0070_em-eta10-phi3*/	2,55,2,11,56,0,1,
/* out0071_em-eta11-phi3*/	6,44,0,1,44,1,10,55,2,1,111,1,2,112,0,14,112,1,4,
/* out0072_em-eta12-phi3*/	6,44,0,4,44,1,1,44,2,4,105,1,4,112,0,2,112,2,9,
/* out0073_em-eta13-phi3*/	7,32,2,1,33,0,1,33,1,2,44,0,1,44,2,3,105,1,8,106,0,3,
/* out0074_em-eta14-phi3*/	6,33,0,6,97,0,3,97,1,2,105,2,2,106,0,1,106,2,1,
/* out0075_em-eta15-phi3*/	4,22,1,1,33,0,4,97,0,2,97,1,5,
/* out0076_em-eta16-phi3*/	4,22,1,3,22,2,1,97,1,1,97,2,6,
/* out0077_em-eta17-phi3*/	4,22,2,4,89,1,1,89,2,4,97,2,1,
/* out0078_em-eta18-phi3*/	2,22,2,3,89,1,4,
/* out0079_em-eta19-phi3*/	1,89,1,2,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	1,95,1,1,
/* out0085_em-eta5-phi4*/	7,88,0,2,88,1,13,95,1,11,95,2,8,96,0,13,96,1,1,96,2,2,
/* out0086_em-eta6-phi4*/	5,77,1,3,78,1,3,88,0,11,88,1,1,88,2,10,
/* out0087_em-eta7-phi4*/	4,67,1,2,77,2,8,78,0,11,78,1,1,
/* out0088_em-eta8-phi4*/	4,67,0,1,67,1,11,67,2,6,78,0,1,
/* out0089_em-eta9-phi4*/	4,56,0,1,56,1,6,67,0,1,67,2,8,
/* out0090_em-eta10-phi4*/	3,56,0,10,56,1,2,56,2,1,
/* out0091_em-eta11-phi4*/	6,44,1,4,44,2,1,45,0,1,56,0,4,56,2,1,112,1,8,
/* out0092_em-eta12-phi4*/	5,44,2,7,45,0,2,106,0,3,112,1,4,112,2,7,
/* out0093_em-eta13-phi4*/	5,33,1,6,44,2,1,106,0,9,106,1,1,106,2,1,
/* out0094_em-eta14-phi4*/	5,33,0,2,33,1,4,33,2,2,97,1,1,106,2,8,
/* out0095_em-eta15-phi4*/	5,33,0,2,33,2,3,97,1,5,98,0,2,106,2,1,
/* out0096_em-eta16-phi4*/	8,23,1,1,23,2,1,33,0,1,33,2,1,97,1,2,97,2,1,98,0,2,98,2,1,
/* out0097_em-eta17-phi4*/	2,23,1,3,89,2,6,
/* out0098_em-eta18-phi4*/	4,23,1,2,89,0,2,89,1,2,89,2,2,
/* out0099_em-eta19-phi4*/	1,89,1,2,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	0,
/* out0105_em-eta5-phi5*/	7,88,1,2,88,2,1,89,0,1,89,1,7,96,0,3,96,1,15,96,2,14,
/* out0106_em-eta6-phi5*/	4,78,1,6,88,2,5,89,0,15,89,1,1,
/* out0107_em-eta7-phi5*/	3,78,0,3,78,1,6,78,2,14,
/* out0108_em-eta8-phi5*/	5,67,2,1,68,0,7,68,1,8,78,0,1,78,2,2,
/* out0109_em-eta9-phi5*/	3,56,1,6,67,2,1,68,0,9,
/* out0110_em-eta10-phi5*/	2,56,1,2,56,2,10,
/* out0111_em-eta11-phi5*/	4,45,1,7,56,2,4,113,0,7,113,1,4,
/* out0112_em-eta12-phi5*/	5,45,0,8,45,1,1,106,1,2,113,0,9,113,2,8,
/* out0113_em-eta13-phi5*/	4,33,1,3,45,0,5,106,1,11,113,2,1,
/* out0114_em-eta14-phi5*/	5,33,1,1,33,2,5,98,0,2,106,1,2,106,2,5,
/* out0115_em-eta15-phi5*/	2,33,2,5,98,0,8,
/* out0116_em-eta16-phi5*/	3,23,2,5,98,0,2,98,2,4,
/* out0117_em-eta17-phi5*/	4,23,1,3,23,2,1,89,2,3,98,2,3,
/* out0118_em-eta18-phi5*/	3,23,1,3,89,0,10,89,2,1,
/* out0119_em-eta19-phi5*/	2,89,0,4,89,1,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	0,
/* out0125_em-eta5-phi6*/	7,89,1,7,89,2,1,90,0,1,90,1,2,97,0,16,97,1,11,97,2,14,
/* out0126_em-eta6-phi6*/	4,79,1,6,89,1,1,89,2,15,90,0,5,
/* out0127_em-eta7-phi6*/	3,79,0,14,79,1,6,79,2,3,
/* out0128_em-eta8-phi6*/	5,68,1,8,68,2,7,69,0,1,79,0,2,79,2,1,
/* out0129_em-eta9-phi6*/	3,57,1,6,68,2,9,69,0,1,
/* out0130_em-eta10-phi6*/	2,57,0,10,57,1,2,
/* out0131_em-eta11-phi6*/	4,45,1,7,57,0,4,113,1,7,114,0,1,
/* out0132_em-eta12-phi6*/	5,45,1,1,45,2,8,107,0,2,113,1,5,113,2,7,
/* out0133_em-eta13-phi6*/	3,34,1,3,45,2,5,107,0,11,
/* out0134_em-eta14-phi6*/	5,34,0,5,34,1,1,98,1,2,107,0,2,107,2,5,
/* out0135_em-eta15-phi6*/	2,34,0,5,98,1,8,
/* out0136_em-eta16-phi6*/	3,23,2,5,98,1,2,98,2,4,
/* out0137_em-eta17-phi6*/	5,23,0,3,23,1,1,23,2,2,90,2,3,98,2,3,
/* out0138_em-eta18-phi6*/	2,23,1,2,90,1,4,
/* out0139_em-eta19-phi6*/	1,90,1,3,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	1,98,1,1,
/* out0145_em-eta5-phi7*/	7,90,1,13,90,2,2,97,1,5,97,2,2,98,0,16,98,1,6,98,2,8,
/* out0146_em-eta6-phi7*/	5,79,1,3,80,1,3,90,0,10,90,1,1,90,2,11,
/* out0147_em-eta7-phi7*/	4,69,1,2,79,1,1,79,2,11,80,0,8,
/* out0148_em-eta8-phi7*/	4,69,0,6,69,1,11,69,2,1,79,2,1,
/* out0149_em-eta9-phi7*/	4,57,1,6,57,2,1,69,0,8,69,2,1,
/* out0150_em-eta10-phi7*/	3,57,0,1,57,1,2,57,2,10,
/* out0151_em-eta11-phi7*/	7,45,2,1,46,0,1,46,1,4,57,0,1,57,2,4,114,0,8,114,1,6,
/* out0152_em-eta12-phi7*/	5,45,2,2,46,0,7,107,1,3,114,0,7,114,2,7,
/* out0153_em-eta13-phi7*/	5,34,1,6,46,0,1,107,0,1,107,1,9,107,2,1,
/* out0154_em-eta14-phi7*/	5,34,0,2,34,1,4,34,2,2,99,0,1,107,2,8,
/* out0155_em-eta15-phi7*/	5,34,0,3,34,2,2,98,1,2,99,0,5,107,2,1,
/* out0156_em-eta16-phi7*/	8,23,0,2,23,2,2,34,0,1,34,2,1,98,1,2,98,2,1,99,0,2,99,2,1,
/* out0157_em-eta17-phi7*/	2,23,0,8,90,2,6,
/* out0158_em-eta18-phi7*/	4,23,0,3,23,1,1,90,1,2,90,2,2,
/* out0159_em-eta19-phi7*/	1,90,1,3,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	1,98,1,3,
/* out0165_em-eta5-phi8*/	9,90,2,1,91,0,5,91,1,14,91,2,1,98,1,6,98,2,8,99,0,4,99,1,3,99,2,1,
/* out0166_em-eta6-phi8*/	5,80,1,11,80,2,2,90,2,2,91,0,11,91,2,2,
/* out0167_em-eta7-phi8*/	4,70,1,1,80,0,8,80,1,2,80,2,12,
/* out0168_em-eta8-phi8*/	4,69,1,3,69,2,9,70,0,5,70,1,1,
/* out0169_em-eta9-phi8*/	3,58,0,1,58,1,9,69,2,5,
/* out0170_em-eta10-phi8*/	2,57,2,1,58,0,11,
/* out0171_em-eta11-phi8*/	5,46,1,10,46,2,1,58,0,1,114,1,9,115,0,2,
/* out0172_em-eta12-phi8*/	6,46,0,4,46,1,1,46,2,4,108,0,4,114,1,1,114,2,9,
/* out0173_em-eta13-phi8*/	7,34,1,2,34,2,1,35,0,1,46,0,3,46,2,1,107,1,3,108,0,8,
/* out0174_em-eta14-phi8*/	6,34,2,6,99,0,2,99,1,3,107,1,1,107,2,1,108,2,2,
/* out0175_em-eta15-phi8*/	4,24,1,1,34,2,4,99,0,5,99,1,2,
/* out0176_em-eta16-phi8*/	4,24,0,1,24,1,3,99,0,1,99,2,6,
/* out0177_em-eta17-phi8*/	4,24,0,4,90,0,1,90,2,4,99,2,1,
/* out0178_em-eta18-phi8*/	4,24,0,3,90,0,6,90,1,1,90,2,1,
/* out0179_em-eta19-phi8*/	1,90,1,2,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	4,92,1,1,99,0,2,99,1,1,99,2,4,
/* out0185_em-eta5-phi9*/	7,91,1,2,91,2,7,92,0,10,92,1,8,99,0,10,99,1,12,99,2,11,
/* out0186_em-eta6-phi9*/	5,81,0,6,81,1,14,81,2,1,91,2,6,92,0,1,
/* out0187_em-eta7-phi9*/	5,70,1,10,70,2,1,80,2,2,81,0,10,81,2,1,
/* out0188_em-eta8-phi9*/	3,70,0,8,70,1,4,70,2,7,
/* out0189_em-eta9-phi9*/	5,58,1,7,58,2,5,59,0,1,70,0,3,70,2,1,
/* out0190_em-eta10-phi9*/	3,47,1,1,58,0,2,58,2,10,
/* out0191_em-eta11-phi9*/	7,46,1,1,46,2,3,47,0,3,47,1,2,58,0,1,115,0,11,115,2,3,
/* out0192_em-eta12-phi9*/	7,35,1,2,46,2,6,47,0,1,108,0,2,108,1,7,115,0,1,115,2,5,
/* out0193_em-eta13-phi9*/	6,35,0,2,35,1,5,46,2,1,108,0,2,108,1,3,108,2,5,
/* out0194_em-eta14-phi9*/	4,35,0,6,99,1,3,100,0,1,108,2,5,
/* out0195_em-eta15-phi9*/	4,24,1,4,35,0,1,99,1,7,99,2,1,
/* out0196_em-eta16-phi9*/	3,24,1,4,91,0,1,99,2,6,
/* out0197_em-eta17-phi9*/	4,24,0,3,90,0,2,91,0,3,99,2,1,
/* out0198_em-eta18-phi9*/	3,24,0,3,90,0,6,91,0,2,
/* out0199_em-eta19-phi9*/	2,90,0,1,90,1,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	2,92,1,2,93,0,1,
/* out0205_em-eta5-phi10*/	6,82,1,4,92,0,3,92,1,5,92,2,15,93,0,8,93,2,1,
/* out0206_em-eta6-phi10*/	6,81,1,2,81,2,9,82,0,9,82,1,4,92,0,2,92,2,1,
/* out0207_em-eta7-phi10*/	4,70,2,1,71,0,5,71,1,10,81,2,5,
/* out0208_em-eta8-phi10*/	3,59,1,6,70,2,6,71,0,6,
/* out0209_em-eta9-phi10*/	2,59,0,9,59,1,6,
/* out0210_em-eta10-phi10*/	3,47,1,8,58,2,1,59,0,4,
/* out0211_em-eta11-phi10*/	6,47,0,5,47,1,4,47,2,2,109,0,2,115,0,2,115,2,5,
/* out0212_em-eta12-phi10*/	5,35,1,3,47,0,6,108,1,3,109,0,9,115,2,3,
/* out0213_em-eta13-phi10*/	8,35,1,5,35,2,2,100,0,1,100,1,1,108,1,3,108,2,3,109,0,2,109,2,1,
/* out0214_em-eta14-phi10*/	4,35,0,4,35,2,3,100,0,8,108,2,1,
/* out0215_em-eta15-phi10*/	5,24,1,3,35,0,2,99,1,1,100,0,5,100,2,2,
/* out0216_em-eta16-phi10*/	4,24,1,1,24,2,3,91,0,3,91,1,3,
/* out0217_em-eta17-phi10*/	2,24,2,4,91,0,5,
/* out0218_em-eta18-phi10*/	4,24,0,1,24,2,2,91,0,2,91,2,3,
/* out0219_em-eta19-phi10*/	2,24,0,1,91,2,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	0,
/* out0225_em-eta5-phi11*/	6,82,1,6,82,2,2,83,0,3,83,1,4,93,0,7,93,2,15,
/* out0226_em-eta6-phi11*/	5,72,1,4,82,0,7,82,1,2,82,2,14,83,0,1,
/* out0227_em-eta7-phi11*/	4,71,0,1,71,1,6,71,2,12,72,0,4,
/* out0228_em-eta8-phi11*/	6,59,1,3,59,2,2,60,0,3,60,1,4,71,0,4,71,2,4,
/* out0229_em-eta9-phi11*/	4,48,1,1,59,1,1,59,2,12,60,0,1,
/* out0230_em-eta10-phi11*/	6,47,1,1,47,2,2,48,0,3,48,1,3,59,0,2,59,2,2,
/* out0231_em-eta11-phi11*/	4,36,1,1,47,2,9,48,0,1,109,1,6,
/* out0232_em-eta12-phi11*/	8,35,1,1,36,0,2,36,1,3,47,0,1,47,2,3,109,0,3,109,1,6,109,2,4,
/* out0233_em-eta13-phi11*/	4,35,2,5,36,0,2,100,1,4,109,2,7,
/* out0234_em-eta14-phi11*/	5,25,1,2,35,2,5,100,0,1,100,1,7,100,2,1,
/* out0235_em-eta15-phi11*/	4,25,0,2,25,1,2,35,2,1,100,2,8,
/* out0236_em-eta16-phi11*/	4,24,2,3,25,0,2,91,1,5,100,2,1,
/* out0237_em-eta17-phi11*/	4,14,1,1,24,2,3,91,1,4,91,2,2,
/* out0238_em-eta18-phi11*/	3,14,1,3,24,2,1,91,2,5,
/* out0239_em-eta19-phi11*/	2,14,1,1,91,2,2,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	0,
/* out0245_em-eta5-phi12*/	4,83,0,6,83,1,12,83,2,13,84,0,3,
/* out0246_em-eta6-phi12*/	6,72,1,12,72,2,6,73,0,1,73,1,1,83,0,6,83,2,1,
/* out0247_em-eta7-phi12*/	4,60,1,4,60,2,1,72,0,12,72,2,6,
/* out0248_em-eta8-phi12*/	3,60,0,5,60,1,8,60,2,6,
/* out0249_em-eta9-phi12*/	3,48,1,8,60,0,7,60,2,1,
/* out0250_em-eta10-phi12*/	3,48,0,5,48,1,4,48,2,3,
/* out0251_em-eta11-phi12*/	4,36,1,5,48,0,6,109,1,1,110,0,8,
/* out0252_em-eta12-phi12*/	9,36,0,2,36,1,6,36,2,1,101,0,2,101,1,2,109,1,3,109,2,3,110,0,4,110,2,2,
/* out0253_em-eta13-phi12*/	3,36,0,8,101,0,9,109,2,1,
/* out0254_em-eta14-phi12*/	5,25,1,6,92,1,1,100,1,4,100,2,1,101,0,3,
/* out0255_em-eta15-phi12*/	4,25,0,2,25,1,3,92,0,5,100,2,3,
/* out0256_em-eta16-phi12*/	3,25,0,5,91,1,1,92,0,5,
/* out0257_em-eta17-phi12*/	6,14,1,1,14,2,2,25,0,1,91,1,3,91,2,1,92,0,1,
/* out0258_em-eta18-phi12*/	3,14,1,4,83,1,3,91,2,2,
/* out0259_em-eta19-phi12*/	2,14,1,1,83,1,2,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	1,84,0,3,
/* out0265_em-eta5-phi13*/	6,73,1,10,73,2,3,74,0,1,83,2,2,84,0,10,84,2,14,
/* out0266_em-eta6-phi13*/	5,61,1,2,72,2,2,73,0,15,73,1,5,73,2,4,
/* out0267_em-eta7-phi13*/	4,61,0,6,61,1,13,61,2,1,72,2,2,
/* out0268_em-eta8-phi13*/	3,49,1,6,60,2,7,61,0,6,
/* out0269_em-eta9-phi13*/	4,48,2,3,49,0,7,49,1,5,60,2,1,
/* out0270_em-eta10-phi13*/	3,37,1,3,48,2,9,49,0,1,
/* out0271_em-eta11-phi13*/	8,36,1,1,36,2,2,37,0,3,37,1,3,48,0,1,48,2,1,110,0,4,110,2,6,
/* out0272_em-eta12-phi13*/	4,36,2,9,101,1,6,102,0,1,110,2,7,
/* out0273_em-eta13-phi13*/	6,26,1,1,36,0,2,36,2,4,101,0,2,101,1,5,101,2,4,
/* out0274_em-eta14-phi13*/	4,25,1,3,25,2,3,92,1,2,101,2,7,
/* out0275_em-eta15-phi13*/	3,25,2,5,92,0,2,92,1,6,
/* out0276_em-eta16-phi13*/	4,25,0,3,25,2,1,92,0,3,92,2,4,
/* out0277_em-eta17-phi13*/	4,14,2,4,25,0,1,83,2,3,92,2,3,
/* out0278_em-eta18-phi13*/	4,14,1,2,14,2,3,83,1,5,83,2,1,
/* out0279_em-eta19-phi13*/	2,14,1,1,83,1,2,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	3,74,0,1,74,1,1,84,2,1,
/* out0285_em-eta5-phi14*/	5,73,2,2,74,0,14,74,1,9,74,2,15,84,2,1,
/* out0286_em-eta6-phi14*/	5,61,1,1,61,2,1,62,0,5,62,1,13,73,2,7,
/* out0287_em-eta7-phi14*/	4,50,1,4,61,0,1,61,2,13,62,0,5,
/* out0288_em-eta8-phi14*/	6,49,1,4,49,2,5,50,0,3,50,1,2,61,0,3,61,2,1,
/* out0289_em-eta9-phi14*/	3,49,0,6,49,1,1,49,2,9,
/* out0290_em-eta10-phi14*/	3,37,1,8,37,2,2,49,0,2,
/* out0291_em-eta11-phi14*/	6,37,0,7,37,1,2,37,2,2,102,0,4,102,1,6,110,2,1,
/* out0292_em-eta12-phi14*/	5,26,1,5,37,0,4,101,1,1,102,0,10,102,2,2,
/* out0293_em-eta13-phi14*/	8,26,0,2,26,1,6,93,0,3,93,1,1,101,1,2,101,2,3,102,0,1,102,2,1,
/* out0294_em-eta14-phi14*/	5,25,2,1,26,0,5,92,1,1,93,0,6,101,2,2,
/* out0295_em-eta15-phi14*/	6,15,1,1,25,2,4,26,0,1,92,1,6,92,2,1,93,0,1,
/* out0296_em-eta16-phi14*/	3,15,1,3,25,2,2,92,2,6,
/* out0297_em-eta17-phi14*/	5,14,2,3,15,0,2,83,2,4,84,0,1,92,2,2,
/* out0298_em-eta18-phi14*/	4,14,1,1,14,2,3,83,1,2,83,2,4,
/* out0299_em-eta19-phi14*/	2,14,1,1,83,1,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	0,
/* out0305_em-eta5-phi15*/	5,62,1,1,63,0,5,63,1,15,74,1,6,74,2,1,
/* out0306_em-eta6-phi15*/	5,51,1,4,62,0,2,62,1,2,62,2,15,63,0,5,
/* out0307_em-eta7-phi15*/	6,50,1,9,50,2,7,51,0,2,51,1,1,62,0,4,62,2,1,
/* out0308_em-eta8-phi15*/	4,38,1,1,50,0,13,50,1,1,50,2,3,
/* out0309_em-eta9-phi15*/	3,38,0,1,38,1,13,49,2,2,
/* out0310_em-eta10-phi15*/	2,37,2,5,38,0,8,
/* out0311_em-eta11-phi15*/	8,27,1,3,37,0,1,37,2,7,102,1,9,102,2,1,103,0,10,103,1,7,103,2,3,
/* out0312_em-eta12-phi15*/	8,26,1,3,26,2,3,27,0,1,27,1,1,37,0,1,94,0,1,102,1,1,102,2,11,
/* out0313_em-eta13-phi15*/	5,26,0,1,26,1,1,26,2,5,93,1,9,102,2,1,
/* out0314_em-eta14-phi15*/	4,26,0,6,93,0,4,93,1,2,93,2,4,
/* out0315_em-eta15-phi15*/	4,15,1,5,84,1,2,93,0,2,93,2,3,
/* out0316_em-eta16-phi15*/	4,15,0,1,15,1,3,84,0,5,84,1,1,
/* out0317_em-eta17-phi15*/	3,15,0,4,83,2,1,84,0,5,
/* out0318_em-eta18-phi15*/	5,14,2,1,15,0,1,83,1,1,83,2,3,84,0,1,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	2,64,0,1,64,2,1,
/* out0325_em-eta5-phi16*/	7,52,1,8,63,0,2,63,1,1,63,2,16,64,0,14,64,1,13,64,2,11,
/* out0326_em-eta6-phi16*/	4,51,1,11,51,2,9,52,0,3,63,0,4,
/* out0327_em-eta7-phi16*/	4,39,1,5,50,2,3,51,0,13,51,2,1,
/* out0328_em-eta8-phi16*/	5,38,1,1,38,2,1,39,0,5,39,1,8,50,2,3,
/* out0329_em-eta9-phi16*/	4,38,0,1,38,1,1,38,2,13,39,0,1,
/* out0330_em-eta10-phi16*/	4,27,1,4,27,2,1,38,0,6,38,2,2,
/* out0331_em-eta11-phi16*/	7,27,0,2,27,1,8,27,2,1,94,1,5,103,0,6,103,1,9,103,2,13,
/* out0332_em-eta12-phi16*/	4,26,2,1,27,0,8,94,0,10,94,1,3,
/* out0333_em-eta13-phi16*/	5,16,1,3,26,2,5,93,1,4,94,0,5,94,2,1,
/* out0334_em-eta14-phi16*/	8,15,1,1,15,2,1,16,0,1,16,1,2,26,0,1,26,2,2,85,0,2,93,2,7,
/* out0335_em-eta15-phi16*/	5,15,1,2,15,2,3,84,1,5,85,0,1,93,2,2,
/* out0336_em-eta16-phi16*/	6,15,0,1,15,1,1,15,2,3,84,0,1,84,1,4,84,2,1,
/* out0337_em-eta17-phi16*/	3,15,0,4,84,0,2,84,2,3,
/* out0338_em-eta18-phi16*/	3,15,0,1,84,0,1,84,2,2,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	0,
/* out0345_em-eta5-phi17*/	9,52,0,2,52,1,8,52,2,15,53,0,12,53,1,8,53,2,4,64,0,1,64,1,3,64,2,4,
/* out0346_em-eta6-phi17*/	4,40,1,12,51,2,4,52,0,11,52,2,1,
/* out0347_em-eta7-phi17*/	6,39,1,2,39,2,6,40,0,8,40,1,4,51,0,1,51,2,2,
/* out0348_em-eta8-phi17*/	3,39,0,8,39,1,1,39,2,10,
/* out0349_em-eta9-phi17*/	2,28,1,13,39,0,2,
/* out0350_em-eta10-phi17*/	3,27,2,3,28,0,8,28,1,3,
/* out0351_em-eta11-phi17*/	5,27,2,10,94,1,4,95,0,12,95,1,8,95,2,4,
/* out0352_em-eta12-phi17*/	5,16,1,3,27,0,5,27,2,1,94,1,4,94,2,9,
/* out0353_em-eta13-phi17*/	3,16,1,7,85,1,6,94,2,6,
/* out0354_em-eta14-phi17*/	4,16,0,5,16,1,1,85,0,7,85,1,2,
/* out0355_em-eta15-phi17*/	4,15,2,3,16,0,2,84,1,2,85,0,6,
/* out0356_em-eta16-phi17*/	3,15,2,4,84,1,2,84,2,4,
/* out0357_em-eta17-phi17*/	3,15,0,2,15,2,2,84,2,5,
/* out0358_em-eta18-phi17*/	1,84,2,1,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	0,
/* out0365_em-eta5-phi18*/	9,41,0,2,41,1,15,41,2,8,42,0,4,42,1,3,42,2,1,53,0,4,53,1,8,53,2,12,
/* out0366_em-eta6-phi18*/	4,30,1,4,40,2,12,41,0,11,41,1,1,
/* out0367_em-eta7-phi18*/	6,29,1,6,29,2,2,30,0,1,30,1,2,40,0,8,40,2,4,
/* out0368_em-eta8-phi18*/	3,29,0,8,29,1,10,29,2,1,
/* out0369_em-eta9-phi18*/	2,28,2,13,29,0,2,
/* out0370_em-eta10-phi18*/	3,17,1,3,28,0,8,28,2,3,
/* out0371_em-eta11-phi18*/	5,17,1,10,86,1,4,95,0,4,95,1,8,95,2,12,
/* out0372_em-eta12-phi18*/	5,16,2,3,17,0,5,17,1,1,86,0,9,86,1,4,
/* out0373_em-eta13-phi18*/	3,16,2,7,85,1,6,86,0,6,
/* out0374_em-eta14-phi18*/	4,16,0,5,16,2,1,85,1,2,85,2,7,
/* out0375_em-eta15-phi18*/	4,7,1,3,16,0,2,80,1,2,85,2,6,
/* out0376_em-eta16-phi18*/	3,7,1,4,80,0,4,80,1,2,
/* out0377_em-eta17-phi18*/	3,7,0,2,7,1,2,80,0,5,
/* out0378_em-eta18-phi18*/	1,80,0,1,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	2,42,0,1,42,2,1,
/* out0385_em-eta5-phi19*/	7,31,0,2,31,1,16,31,2,1,41,2,8,42,0,11,42,1,13,42,2,14,
/* out0386_em-eta6-phi19*/	4,30,1,9,30,2,11,31,0,4,41,0,3,
/* out0387_em-eta7-phi19*/	4,19,1,3,29,2,5,30,0,13,30,1,1,
/* out0388_em-eta8-phi19*/	5,18,1,1,18,2,1,19,1,3,29,0,5,29,2,8,
/* out0389_em-eta9-phi19*/	4,18,0,1,18,1,13,18,2,1,29,0,1,
/* out0390_em-eta10-phi19*/	4,17,1,1,17,2,4,18,0,6,18,1,2,
/* out0391_em-eta11-phi19*/	7,17,0,2,17,1,1,17,2,8,86,1,5,87,0,13,87,1,9,87,2,6,
/* out0392_em-eta12-phi19*/	4,8,1,1,17,0,8,86,1,3,86,2,10,
/* out0393_em-eta13-phi19*/	5,8,1,5,16,2,3,81,1,4,86,0,1,86,2,5,
/* out0394_em-eta14-phi19*/	8,7,1,1,7,2,1,8,0,1,8,1,2,16,0,1,16,2,2,81,0,7,85,2,2,
/* out0395_em-eta15-phi19*/	5,7,1,3,7,2,2,80,1,5,81,0,2,85,2,1,
/* out0396_em-eta16-phi19*/	6,7,0,1,7,1,3,7,2,1,80,0,1,80,1,4,80,2,1,
/* out0397_em-eta17-phi19*/	3,7,0,4,80,0,3,80,2,2,
/* out0398_em-eta18-phi19*/	3,7,0,1,80,0,2,80,2,1,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	0,
/* out0405_em-eta5-phi20*/	6,20,2,1,21,0,13,21,1,2,21,2,1,31,0,5,31,2,15,
/* out0406_em-eta6-phi20*/	5,20,0,2,20,1,15,20,2,2,30,2,4,31,0,5,
/* out0407_em-eta7-phi20*/	6,19,1,7,19,2,9,20,0,4,20,1,1,30,0,2,30,2,1,
/* out0408_em-eta8-phi20*/	4,18,2,1,19,0,13,19,1,3,19,2,1,
/* out0409_em-eta9-phi20*/	3,10,1,2,18,0,1,18,2,13,
/* out0410_em-eta10-phi20*/	2,9,1,5,18,0,8,
/* out0411_em-eta11-phi20*/	8,9,0,1,9,1,7,17,2,3,82,0,1,82,1,9,87,0,3,87,1,7,87,2,10,
/* out0412_em-eta12-phi20*/	8,8,1,3,8,2,3,9,0,1,17,0,1,17,2,1,82,0,11,82,1,1,86,2,1,
/* out0413_em-eta13-phi20*/	5,8,0,1,8,1,5,8,2,1,81,1,9,82,0,1,
/* out0414_em-eta14-phi20*/	4,8,0,6,81,0,4,81,1,2,81,2,4,
/* out0415_em-eta15-phi20*/	4,7,2,5,80,1,2,81,0,3,81,2,2,
/* out0416_em-eta16-phi20*/	4,7,0,1,7,2,3,80,1,1,80,2,5,
/* out0417_em-eta17-phi20*/	3,7,0,4,76,1,1,80,2,5,
/* out0418_em-eta18-phi20*/	4,0,1,2,7,0,1,76,1,4,80,2,1,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	2,13,0,1,21,1,1,
/* out0425_em-eta5-phi21*/	5,12,1,2,13,0,1,21,0,3,21,1,13,21,2,15,
/* out0426_em-eta6-phi21*/	5,11,1,1,11,2,1,12,1,7,20,0,5,20,2,13,
/* out0427_em-eta7-phi21*/	4,11,0,1,11,1,13,19,2,4,20,0,5,
/* out0428_em-eta8-phi21*/	6,10,1,5,10,2,4,11,0,3,11,1,1,19,0,3,19,2,2,
/* out0429_em-eta9-phi21*/	3,10,0,6,10,1,9,10,2,1,
/* out0430_em-eta10-phi21*/	3,9,1,2,9,2,8,10,0,2,
/* out0431_em-eta11-phi21*/	6,9,0,7,9,1,2,9,2,2,79,0,1,82,1,6,82,2,4,
/* out0432_em-eta12-phi21*/	5,8,2,5,9,0,4,78,1,1,82,0,2,82,2,10,
/* out0433_em-eta13-phi21*/	8,8,0,2,8,2,6,78,0,3,78,1,2,81,1,1,81,2,3,82,0,1,82,2,1,
/* out0434_em-eta14-phi21*/	5,1,1,1,8,0,5,77,1,1,78,0,2,81,2,6,
/* out0435_em-eta15-phi21*/	6,1,1,4,7,2,1,8,0,1,77,0,1,77,1,6,81,2,1,
/* out0436_em-eta16-phi21*/	3,1,1,2,7,2,3,77,0,6,
/* out0437_em-eta17-phi21*/	8,0,1,3,0,2,1,1,0,1,7,0,2,76,1,1,76,2,2,77,0,2,80,2,1,
/* out0438_em-eta18-phi21*/	3,0,1,4,76,1,5,76,2,1,
/* out0439_em-eta19-phi21*/	1,76,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	1,13,0,3,
/* out0445_em-eta5-phi22*/	5,6,1,2,12,1,3,12,2,10,13,0,10,13,2,14,
/* out0446_em-eta6-phi22*/	5,5,1,2,11,2,2,12,0,15,12,1,4,12,2,5,
/* out0447_em-eta7-phi22*/	4,5,1,2,11,0,6,11,1,1,11,2,13,
/* out0448_em-eta8-phi22*/	3,4,1,7,10,2,6,11,0,6,
/* out0449_em-eta9-phi22*/	6,3,1,3,3,2,3,4,0,3,4,1,1,10,0,7,10,2,5,
/* out0450_em-eta10-phi22*/	3,3,1,9,9,2,3,10,0,1,
/* out0451_em-eta11-phi22*/	8,2,1,2,2,2,2,3,0,1,3,1,1,9,0,3,9,2,3,79,0,9,79,2,1,
/* out0452_em-eta12-phi22*/	6,2,1,9,2,2,2,78,1,6,79,0,3,79,2,5,82,2,1,
/* out0453_em-eta13-phi22*/	7,1,2,1,2,0,3,2,1,4,8,2,1,78,0,4,78,1,5,78,2,2,
/* out0454_em-eta14-phi22*/	5,1,1,3,1,2,3,2,0,1,77,1,2,78,0,7,
/* out0455_em-eta15-phi22*/	5,1,0,1,1,1,5,1,2,1,77,1,6,77,2,2,
/* out0456_em-eta16-phi22*/	4,1,0,3,1,1,1,77,0,4,77,2,3,
/* out0457_em-eta17-phi22*/	5,0,1,1,0,2,4,1,0,1,76,2,3,77,0,3,
/* out0458_em-eta18-phi22*/	4,0,1,3,0,2,2,76,1,1,76,2,6,
/* out0459_em-eta19-phi22*/	2,0,1,1,76,1,2,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	0,
/* out0465_em-eta5-phi23*/	5,6,0,6,6,1,13,6,2,16,13,0,1,13,2,2,
/* out0466_em-eta6-phi23*/	6,5,1,6,5,2,12,6,0,10,6,1,1,12,0,1,12,2,1,
/* out0467_em-eta7-phi23*/	5,4,1,1,4,2,8,5,0,16,5,1,6,5,2,4,
/* out0468_em-eta8-phi23*/	3,4,0,5,4,1,6,4,2,8,
/* out0469_em-eta9-phi23*/	3,3,2,8,4,0,8,4,1,1,
/* out0470_em-eta10-phi23*/	3,3,0,9,3,1,3,3,2,5,
/* out0471_em-eta11-phi23*/	4,2,2,6,3,0,6,79,0,3,79,2,4,
/* out0472_em-eta12-phi23*/	6,2,0,3,2,1,1,2,2,6,78,1,2,78,2,2,79,2,6,
/* out0473_em-eta13-phi23*/	2,2,0,8,78,2,9,
/* out0474_em-eta14-phi23*/	4,1,2,8,2,0,1,77,1,1,78,2,3,
/* out0475_em-eta15-phi23*/	3,1,0,3,1,2,3,77,2,5,
/* out0476_em-eta16-phi23*/	2,1,0,5,77,2,5,
/* out0477_em-eta17-phi23*/	3,0,2,4,1,0,2,77,2,1,
/* out0478_em-eta18-phi23*/	3,0,1,1,0,2,4,76,2,3,
/* out0479_em-eta19-phi23*/	4,0,1,1,0,2,1,76,1,1,76,2,1
};