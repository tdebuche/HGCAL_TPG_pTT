parameter integer matrixH [0:4859] = {
/* num inputs = 152(in0-in151) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1433 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	0, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	0, 
/* out0033_had-eta13-phi1*/	0, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	0, 
/* out0036_had-eta16-phi1*/	0, 
/* out0037_had-eta17-phi1*/	0, 
/* out0038_had-eta18-phi1*/	0, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	0, 
/* out0045_had-eta5-phi2*/	0, 
/* out0046_had-eta6-phi2*/	0, 
/* out0047_had-eta7-phi2*/	0, 
/* out0048_had-eta8-phi2*/	0, 
/* out0049_had-eta9-phi2*/	2, 47, 1, 1, 47, 2, 4, 
/* out0050_had-eta10-phi2*/	1, 47, 1, 3, 
/* out0051_had-eta11-phi2*/	2, 46, 1, 2, 46, 2, 4, 
/* out0052_had-eta12-phi2*/	1, 46, 1, 2, 
/* out0053_had-eta13-phi2*/	1, 45, 2, 4, 
/* out0054_had-eta14-phi2*/	1, 45, 1, 3, 
/* out0055_had-eta15-phi2*/	1, 44, 2, 1, 
/* out0056_had-eta16-phi2*/	2, 44, 1, 1, 44, 2, 3, 
/* out0057_had-eta17-phi2*/	1, 44, 1, 3, 
/* out0058_had-eta18-phi2*/	0, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	1, 107, 0, 2, 
/* out0061_had-eta1-phi3*/	2, 106, 0, 2, 107, 0, 6, 
/* out0062_had-eta2-phi3*/	1, 106, 0, 4, 
/* out0063_had-eta3-phi3*/	2, 105, 0, 3, 106, 0, 2, 
/* out0064_had-eta4-phi3*/	1, 105, 0, 4, 
/* out0065_had-eta5-phi3*/	2, 104, 0, 4, 105, 0, 1, 
/* out0066_had-eta6-phi3*/	1, 104, 0, 4, 
/* out0067_had-eta7-phi3*/	0, 
/* out0068_had-eta8-phi3*/	0, 
/* out0069_had-eta9-phi3*/	4, 47, 0, 5, 47, 1, 2, 47, 2, 12, 99, 1, 12, 
/* out0070_had-eta10-phi3*/	5, 46, 2, 4, 47, 0, 2, 47, 1, 10, 98, 1, 1, 98, 2, 11, 
/* out0071_had-eta11-phi3*/	4, 46, 0, 3, 46, 1, 3, 46, 2, 8, 98, 1, 9, 
/* out0072_had-eta12-phi3*/	3, 45, 2, 2, 46, 1, 8, 97, 2, 8, 
/* out0073_had-eta13-phi3*/	3, 45, 0, 1, 45, 2, 9, 97, 1, 7, 
/* out0074_had-eta14-phi3*/	2, 45, 1, 8, 96, 2, 3, 
/* out0075_had-eta15-phi3*/	4, 44, 2, 5, 45, 1, 2, 96, 1, 3, 96, 2, 3, 
/* out0076_had-eta16-phi3*/	3, 44, 1, 1, 44, 2, 4, 96, 1, 2, 
/* out0077_had-eta17-phi3*/	2, 44, 1, 5, 95, 1, 1, 
/* out0078_had-eta18-phi3*/	2, 44, 1, 2, 95, 1, 2, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	1, 107, 0, 2, 
/* out0081_had-eta1-phi4*/	2, 106, 0, 2, 107, 0, 6, 
/* out0082_had-eta2-phi4*/	1, 106, 0, 4, 
/* out0083_had-eta3-phi4*/	2, 105, 0, 3, 106, 0, 2, 
/* out0084_had-eta4-phi4*/	1, 105, 0, 4, 
/* out0085_had-eta5-phi4*/	2, 104, 0, 4, 105, 0, 1, 
/* out0086_had-eta6-phi4*/	1, 104, 0, 4, 
/* out0087_had-eta7-phi4*/	0, 
/* out0088_had-eta8-phi4*/	1, 43, 1, 1, 
/* out0089_had-eta9-phi4*/	7, 42, 2, 3, 43, 1, 12, 47, 0, 6, 93, 1, 1, 93, 2, 5, 99, 0, 16, 99, 1, 4, 
/* out0090_had-eta10-phi4*/	7, 42, 1, 4, 42, 2, 8, 46, 0, 1, 47, 0, 3, 93, 1, 2, 98, 0, 10, 98, 2, 5, 
/* out0091_had-eta11-phi4*/	8, 41, 2, 2, 42, 1, 4, 46, 0, 9, 91, 2, 1, 97, 0, 1, 97, 2, 2, 98, 0, 5, 98, 1, 6, 
/* out0092_had-eta12-phi4*/	8, 41, 1, 2, 41, 2, 4, 45, 0, 1, 45, 2, 1, 46, 0, 3, 46, 1, 1, 97, 0, 6, 97, 2, 6, 
/* out0093_had-eta13-phi4*/	4, 41, 1, 1, 45, 0, 8, 97, 0, 2, 97, 1, 8, 
/* out0094_had-eta14-phi4*/	5, 40, 2, 1, 45, 0, 6, 45, 1, 2, 96, 2, 8, 97, 1, 1, 
/* out0095_had-eta15-phi4*/	7, 40, 1, 1, 44, 0, 2, 44, 2, 2, 45, 1, 1, 96, 0, 1, 96, 1, 4, 96, 2, 2, 
/* out0096_had-eta16-phi4*/	4, 44, 0, 5, 44, 2, 1, 95, 1, 1, 96, 1, 5, 
/* out0097_had-eta17-phi4*/	3, 44, 0, 2, 44, 1, 2, 95, 1, 5, 
/* out0098_had-eta18-phi4*/	2, 44, 1, 2, 95, 1, 3, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	1, 111, 0, 2, 
/* out0101_had-eta1-phi5*/	2, 110, 0, 2, 111, 0, 6, 
/* out0102_had-eta2-phi5*/	1, 110, 0, 4, 
/* out0103_had-eta3-phi5*/	2, 109, 0, 3, 110, 0, 2, 
/* out0104_had-eta4-phi5*/	1, 109, 0, 4, 
/* out0105_had-eta5-phi5*/	2, 108, 0, 4, 109, 0, 1, 
/* out0106_had-eta6-phi5*/	1, 108, 0, 4, 
/* out0107_had-eta7-phi5*/	0, 
/* out0108_had-eta8-phi5*/	2, 37, 2, 2, 43, 0, 7, 
/* out0109_had-eta9-phi5*/	9, 37, 1, 3, 37, 2, 6, 42, 0, 2, 42, 2, 3, 43, 0, 9, 43, 1, 3, 93, 0, 8, 93, 1, 2, 93, 2, 11, 
/* out0110_had-eta10-phi5*/	7, 42, 0, 11, 42, 1, 3, 42, 2, 2, 91, 2, 5, 93, 0, 1, 93, 1, 11, 98, 0, 1, 
/* out0111_had-eta11-phi5*/	6, 41, 0, 1, 41, 2, 6, 42, 0, 1, 42, 1, 5, 91, 1, 5, 91, 2, 9, 
/* out0112_had-eta12-phi5*/	6, 41, 0, 3, 41, 1, 4, 41, 2, 4, 90, 2, 2, 91, 1, 6, 97, 0, 4, 
/* out0113_had-eta13-phi5*/	5, 40, 2, 3, 41, 1, 7, 90, 1, 1, 90, 2, 6, 97, 0, 3, 
/* out0114_had-eta14-phi5*/	3, 40, 2, 8, 90, 1, 3, 96, 0, 5, 
/* out0115_had-eta15-phi5*/	3, 40, 1, 6, 44, 0, 1, 96, 0, 7, 
/* out0116_had-eta16-phi5*/	7, 39, 2, 1, 40, 1, 1, 44, 0, 4, 95, 0, 1, 95, 1, 1, 96, 0, 2, 96, 1, 2, 
/* out0117_had-eta17-phi5*/	4, 39, 2, 3, 44, 0, 2, 95, 0, 5, 95, 1, 2, 
/* out0118_had-eta18-phi5*/	4, 39, 1, 1, 39, 2, 1, 95, 0, 3, 95, 1, 1, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	1, 111, 0, 2, 
/* out0121_had-eta1-phi6*/	2, 110, 0, 2, 111, 0, 6, 
/* out0122_had-eta2-phi6*/	1, 110, 0, 4, 
/* out0123_had-eta3-phi6*/	2, 109, 0, 3, 110, 0, 2, 
/* out0124_had-eta4-phi6*/	1, 109, 0, 4, 
/* out0125_had-eta5-phi6*/	2, 108, 0, 4, 109, 0, 1, 
/* out0126_had-eta6-phi6*/	1, 108, 0, 4, 
/* out0127_had-eta7-phi6*/	0, 
/* out0128_had-eta8-phi6*/	2, 37, 0, 1, 37, 2, 3, 
/* out0129_had-eta9-phi6*/	5, 37, 0, 8, 37, 1, 10, 37, 2, 5, 93, 0, 5, 94, 2, 6, 
/* out0130_had-eta10-phi6*/	8, 36, 2, 11, 37, 1, 3, 42, 0, 2, 91, 0, 3, 91, 2, 1, 93, 0, 2, 94, 1, 6, 94, 2, 5, 
/* out0131_had-eta11-phi6*/	5, 36, 1, 9, 36, 2, 3, 41, 0, 3, 91, 0, 12, 91, 1, 1, 
/* out0132_had-eta12-phi6*/	7, 35, 2, 3, 41, 0, 8, 90, 0, 2, 90, 2, 4, 91, 0, 1, 91, 1, 4, 92, 2, 1, 
/* out0133_had-eta13-phi6*/	9, 35, 1, 1, 35, 2, 1, 40, 0, 2, 40, 2, 2, 41, 0, 1, 41, 1, 2, 90, 0, 3, 90, 1, 2, 90, 2, 4, 
/* out0134_had-eta14-phi6*/	4, 40, 0, 5, 40, 2, 2, 89, 2, 1, 90, 1, 8, 
/* out0135_had-eta15-phi6*/	4, 40, 0, 1, 40, 1, 6, 89, 2, 6, 96, 0, 1, 
/* out0136_had-eta16-phi6*/	4, 39, 2, 4, 40, 1, 1, 89, 1, 3, 89, 2, 3, 
/* out0137_had-eta17-phi6*/	4, 39, 1, 1, 39, 2, 4, 89, 1, 2, 95, 0, 6, 
/* out0138_had-eta18-phi6*/	2, 39, 1, 5, 95, 0, 1, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	1, 115, 0, 2, 
/* out0141_had-eta1-phi7*/	2, 114, 0, 2, 115, 0, 6, 
/* out0142_had-eta2-phi7*/	1, 114, 0, 4, 
/* out0143_had-eta3-phi7*/	2, 113, 0, 3, 114, 0, 2, 
/* out0144_had-eta4-phi7*/	1, 113, 0, 4, 
/* out0145_had-eta5-phi7*/	2, 112, 0, 4, 113, 0, 1, 
/* out0146_had-eta6-phi7*/	1, 112, 0, 4, 
/* out0147_had-eta7-phi7*/	0, 
/* out0148_had-eta8-phi7*/	0, 
/* out0149_had-eta9-phi7*/	5, 37, 0, 7, 38, 1, 3, 38, 2, 14, 94, 0, 8, 94, 2, 4, 
/* out0150_had-eta10-phi7*/	7, 36, 0, 11, 36, 2, 2, 38, 1, 4, 92, 2, 1, 94, 0, 7, 94, 1, 9, 94, 2, 1, 
/* out0151_had-eta11-phi7*/	5, 35, 2, 1, 36, 0, 5, 36, 1, 7, 92, 2, 13, 94, 1, 1, 
/* out0152_had-eta12-phi7*/	5, 35, 0, 1, 35, 2, 10, 90, 0, 2, 92, 1, 9, 92, 2, 1, 
/* out0153_had-eta13-phi7*/	4, 35, 1, 9, 35, 2, 1, 90, 0, 7, 100, 2, 2, 
/* out0154_had-eta14-phi7*/	8, 29, 2, 2, 35, 1, 1, 40, 0, 5, 89, 0, 1, 89, 2, 2, 90, 0, 2, 90, 1, 2, 100, 2, 1, 
/* out0155_had-eta15-phi7*/	6, 29, 1, 1, 29, 2, 2, 40, 0, 3, 40, 1, 1, 89, 0, 3, 89, 2, 4, 
/* out0156_had-eta16-phi7*/	4, 39, 0, 3, 39, 2, 2, 89, 0, 1, 89, 1, 4, 
/* out0157_had-eta17-phi7*/	4, 39, 0, 3, 39, 1, 1, 39, 2, 1, 89, 1, 4, 
/* out0158_had-eta18-phi7*/	1, 39, 1, 6, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	1, 115, 0, 2, 
/* out0161_had-eta1-phi8*/	2, 114, 0, 2, 115, 0, 6, 
/* out0162_had-eta2-phi8*/	1, 114, 0, 4, 
/* out0163_had-eta3-phi8*/	2, 113, 0, 3, 114, 0, 2, 
/* out0164_had-eta4-phi8*/	1, 113, 0, 4, 
/* out0165_had-eta5-phi8*/	2, 112, 0, 4, 113, 0, 1, 
/* out0166_had-eta6-phi8*/	1, 112, 0, 4, 
/* out0167_had-eta7-phi8*/	0, 
/* out0168_had-eta8-phi8*/	0, 
/* out0169_had-eta9-phi8*/	4, 38, 0, 16, 38, 1, 3, 38, 2, 2, 102, 2, 7, 
/* out0170_had-eta10-phi8*/	6, 31, 2, 9, 38, 1, 6, 92, 0, 1, 94, 0, 1, 102, 1, 6, 102, 2, 9, 
/* out0171_had-eta11-phi8*/	5, 31, 1, 7, 31, 2, 6, 35, 0, 1, 92, 0, 12, 102, 1, 2, 
/* out0172_had-eta12-phi8*/	5, 31, 1, 1, 35, 0, 10, 92, 0, 3, 92, 1, 7, 100, 2, 2, 
/* out0173_had-eta13-phi8*/	4, 29, 2, 1, 35, 0, 4, 35, 1, 5, 100, 2, 10, 
/* out0174_had-eta14-phi8*/	3, 29, 2, 8, 100, 1, 6, 100, 2, 1, 
/* out0175_had-eta15-phi8*/	4, 29, 1, 3, 29, 2, 3, 89, 0, 6, 100, 1, 1, 
/* out0176_had-eta16-phi8*/	4, 29, 1, 3, 39, 0, 2, 89, 0, 5, 89, 1, 1, 
/* out0177_had-eta17-phi8*/	2, 39, 0, 5, 89, 1, 2, 
/* out0178_had-eta18-phi8*/	2, 39, 0, 3, 39, 1, 2, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	1, 119, 0, 2, 
/* out0181_had-eta1-phi9*/	2, 118, 0, 2, 119, 0, 6, 
/* out0182_had-eta2-phi9*/	1, 118, 0, 4, 
/* out0183_had-eta3-phi9*/	2, 117, 0, 3, 118, 0, 2, 
/* out0184_had-eta4-phi9*/	1, 117, 0, 4, 
/* out0185_had-eta5-phi9*/	2, 116, 0, 4, 117, 0, 1, 
/* out0186_had-eta6-phi9*/	1, 116, 0, 4, 
/* out0187_had-eta7-phi9*/	0, 
/* out0188_had-eta8-phi9*/	0, 
/* out0189_had-eta9-phi9*/	4, 33, 0, 2, 33, 1, 3, 33, 2, 16, 102, 0, 7, 
/* out0190_had-eta10-phi9*/	7, 31, 0, 10, 31, 2, 1, 33, 1, 6, 101, 2, 1, 102, 0, 9, 102, 1, 6, 103, 2, 1, 
/* out0191_had-eta11-phi9*/	5, 30, 2, 1, 31, 0, 6, 31, 1, 7, 101, 2, 12, 102, 1, 2, 
/* out0192_had-eta12-phi9*/	5, 30, 2, 10, 31, 1, 1, 100, 0, 2, 101, 1, 7, 101, 2, 3, 
/* out0193_had-eta13-phi9*/	4, 29, 0, 1, 30, 1, 5, 30, 2, 4, 100, 0, 10, 
/* out0194_had-eta14-phi9*/	3, 29, 0, 7, 100, 0, 1, 100, 1, 7, 
/* out0195_had-eta15-phi9*/	4, 29, 0, 3, 29, 1, 4, 85, 2, 6, 100, 1, 1, 
/* out0196_had-eta16-phi9*/	4, 24, 2, 2, 29, 1, 4, 85, 1, 1, 85, 2, 5, 
/* out0197_had-eta17-phi9*/	2, 24, 2, 5, 85, 1, 2, 
/* out0198_had-eta18-phi9*/	2, 24, 1, 2, 24, 2, 3, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	1, 119, 0, 2, 
/* out0201_had-eta1-phi10*/	2, 118, 0, 2, 119, 0, 6, 
/* out0202_had-eta2-phi10*/	1, 118, 0, 4, 
/* out0203_had-eta3-phi10*/	2, 117, 0, 3, 118, 0, 2, 
/* out0204_had-eta4-phi10*/	1, 117, 0, 4, 
/* out0205_had-eta5-phi10*/	2, 116, 0, 4, 117, 0, 1, 
/* out0206_had-eta6-phi10*/	1, 116, 0, 4, 
/* out0207_had-eta7-phi10*/	0, 
/* out0208_had-eta8-phi10*/	0, 
/* out0209_had-eta9-phi10*/	5, 33, 0, 14, 33, 1, 3, 34, 2, 7, 103, 0, 4, 103, 2, 8, 
/* out0210_had-eta10-phi10*/	7, 32, 0, 2, 32, 2, 11, 33, 1, 4, 101, 0, 1, 103, 0, 1, 103, 1, 9, 103, 2, 7, 
/* out0211_had-eta11-phi10*/	5, 30, 0, 1, 32, 1, 7, 32, 2, 5, 101, 0, 13, 103, 1, 1, 
/* out0212_had-eta12-phi10*/	5, 30, 0, 10, 30, 2, 1, 86, 2, 2, 101, 0, 1, 101, 1, 9, 
/* out0213_had-eta13-phi10*/	4, 30, 0, 1, 30, 1, 9, 86, 2, 7, 100, 0, 2, 
/* out0214_had-eta14-phi10*/	9, 25, 2, 5, 29, 0, 2, 30, 1, 1, 85, 0, 2, 85, 2, 1, 86, 1, 2, 86, 2, 2, 100, 0, 1, 100, 1, 1, 
/* out0215_had-eta15-phi10*/	6, 25, 1, 1, 25, 2, 3, 29, 0, 3, 29, 1, 1, 85, 0, 4, 85, 2, 3, 
/* out0216_had-eta16-phi10*/	4, 24, 0, 2, 24, 2, 3, 85, 1, 4, 85, 2, 1, 
/* out0217_had-eta17-phi10*/	4, 24, 0, 1, 24, 1, 1, 24, 2, 3, 85, 1, 4, 
/* out0218_had-eta18-phi10*/	1, 24, 1, 6, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	1, 123, 0, 2, 
/* out0221_had-eta1-phi11*/	2, 122, 0, 2, 123, 0, 6, 
/* out0222_had-eta2-phi11*/	1, 122, 0, 4, 
/* out0223_had-eta3-phi11*/	2, 121, 0, 3, 122, 0, 2, 
/* out0224_had-eta4-phi11*/	1, 121, 0, 4, 
/* out0225_had-eta5-phi11*/	2, 120, 0, 4, 121, 0, 1, 
/* out0226_had-eta6-phi11*/	1, 120, 0, 4, 
/* out0227_had-eta7-phi11*/	0, 
/* out0228_had-eta8-phi11*/	2, 34, 0, 3, 34, 2, 1, 
/* out0229_had-eta9-phi11*/	5, 34, 0, 5, 34, 1, 10, 34, 2, 8, 88, 2, 5, 103, 0, 6, 
/* out0230_had-eta10-phi11*/	8, 27, 2, 2, 32, 0, 11, 34, 1, 3, 87, 0, 1, 87, 2, 3, 88, 2, 2, 103, 0, 5, 103, 1, 6, 
/* out0231_had-eta11-phi11*/	5, 26, 2, 3, 32, 0, 3, 32, 1, 9, 87, 1, 1, 87, 2, 12, 
/* out0232_had-eta12-phi11*/	7, 26, 2, 8, 30, 0, 3, 86, 0, 4, 86, 2, 2, 87, 1, 4, 87, 2, 1, 101, 0, 1, 
/* out0233_had-eta13-phi11*/	9, 25, 0, 2, 25, 2, 2, 26, 1, 2, 26, 2, 1, 30, 0, 1, 30, 1, 1, 86, 0, 4, 86, 1, 2, 86, 2, 3, 
/* out0234_had-eta14-phi11*/	4, 25, 0, 2, 25, 2, 5, 85, 0, 1, 86, 1, 8, 
/* out0235_had-eta15-phi11*/	4, 25, 1, 6, 25, 2, 1, 81, 2, 1, 85, 0, 6, 
/* out0236_had-eta16-phi11*/	4, 24, 0, 4, 25, 1, 1, 85, 0, 3, 85, 1, 3, 
/* out0237_had-eta17-phi11*/	4, 24, 0, 4, 24, 1, 1, 80, 1, 6, 85, 1, 2, 
/* out0238_had-eta18-phi11*/	2, 24, 1, 5, 80, 1, 1, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	1, 123, 0, 2, 
/* out0241_had-eta1-phi12*/	2, 122, 0, 2, 123, 0, 6, 
/* out0242_had-eta2-phi12*/	1, 122, 0, 4, 
/* out0243_had-eta3-phi12*/	2, 121, 0, 3, 122, 0, 2, 
/* out0244_had-eta4-phi12*/	1, 121, 0, 4, 
/* out0245_had-eta5-phi12*/	2, 120, 0, 4, 121, 0, 1, 
/* out0246_had-eta6-phi12*/	1, 120, 0, 4, 
/* out0247_had-eta7-phi12*/	0, 
/* out0248_had-eta8-phi12*/	2, 28, 1, 7, 34, 0, 2, 
/* out0249_had-eta9-phi12*/	9, 27, 0, 3, 27, 2, 2, 28, 0, 3, 28, 1, 9, 34, 0, 6, 34, 1, 3, 88, 0, 11, 88, 1, 2, 88, 2, 8, 
/* out0250_had-eta10-phi12*/	7, 27, 0, 2, 27, 1, 3, 27, 2, 11, 83, 2, 1, 87, 0, 5, 88, 1, 11, 88, 2, 1, 
/* out0251_had-eta11-phi12*/	6, 26, 0, 6, 26, 2, 1, 27, 1, 5, 27, 2, 1, 87, 0, 9, 87, 1, 5, 
/* out0252_had-eta12-phi12*/	6, 26, 0, 4, 26, 1, 4, 26, 2, 3, 82, 2, 4, 86, 0, 2, 87, 1, 6, 
/* out0253_had-eta13-phi12*/	5, 25, 0, 3, 26, 1, 7, 82, 2, 3, 86, 0, 6, 86, 1, 1, 
/* out0254_had-eta14-phi12*/	3, 25, 0, 8, 81, 2, 5, 86, 1, 3, 
/* out0255_had-eta15-phi12*/	3, 20, 2, 1, 25, 1, 6, 81, 2, 7, 
/* out0256_had-eta16-phi12*/	7, 20, 2, 4, 24, 0, 1, 25, 1, 1, 80, 0, 1, 80, 1, 1, 81, 1, 2, 81, 2, 2, 
/* out0257_had-eta17-phi12*/	4, 20, 2, 2, 24, 0, 3, 80, 0, 2, 80, 1, 5, 
/* out0258_had-eta18-phi12*/	4, 24, 0, 1, 24, 1, 1, 80, 0, 1, 80, 1, 3, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	1, 127, 0, 2, 
/* out0261_had-eta1-phi13*/	2, 126, 0, 2, 127, 0, 6, 
/* out0262_had-eta2-phi13*/	1, 126, 0, 4, 
/* out0263_had-eta3-phi13*/	2, 125, 0, 3, 126, 0, 2, 
/* out0264_had-eta4-phi13*/	1, 125, 0, 4, 
/* out0265_had-eta5-phi13*/	2, 124, 0, 4, 125, 0, 1, 
/* out0266_had-eta6-phi13*/	1, 124, 0, 4, 
/* out0267_had-eta7-phi13*/	0, 
/* out0268_had-eta8-phi13*/	1, 28, 0, 1, 
/* out0269_had-eta9-phi13*/	7, 23, 2, 6, 27, 0, 3, 28, 0, 12, 84, 0, 4, 84, 1, 16, 88, 0, 5, 88, 1, 1, 
/* out0270_had-eta10-phi13*/	7, 22, 2, 1, 23, 2, 3, 27, 0, 8, 27, 1, 4, 83, 0, 5, 83, 2, 10, 88, 1, 2, 
/* out0271_had-eta11-phi13*/	8, 22, 2, 9, 26, 0, 2, 27, 1, 4, 82, 0, 2, 82, 2, 1, 83, 1, 6, 83, 2, 5, 87, 0, 1, 
/* out0272_had-eta12-phi13*/	8, 21, 0, 1, 21, 2, 1, 22, 1, 1, 22, 2, 3, 26, 0, 4, 26, 1, 2, 82, 0, 6, 82, 2, 6, 
/* out0273_had-eta13-phi13*/	4, 21, 2, 8, 26, 1, 1, 82, 1, 8, 82, 2, 2, 
/* out0274_had-eta14-phi13*/	5, 21, 1, 2, 21, 2, 6, 25, 0, 1, 81, 0, 8, 82, 1, 1, 
/* out0275_had-eta15-phi13*/	7, 20, 0, 2, 20, 2, 2, 21, 1, 1, 25, 1, 1, 81, 0, 2, 81, 1, 4, 81, 2, 1, 
/* out0276_had-eta16-phi13*/	4, 20, 0, 1, 20, 2, 5, 80, 0, 1, 81, 1, 5, 
/* out0277_had-eta17-phi13*/	3, 20, 1, 2, 20, 2, 2, 80, 0, 5, 
/* out0278_had-eta18-phi13*/	2, 20, 1, 2, 80, 0, 3, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	1, 127, 0, 2, 
/* out0281_had-eta1-phi14*/	2, 126, 0, 2, 127, 0, 6, 
/* out0282_had-eta2-phi14*/	1, 126, 0, 4, 
/* out0283_had-eta3-phi14*/	2, 125, 0, 3, 126, 0, 2, 
/* out0284_had-eta4-phi14*/	1, 125, 0, 4, 
/* out0285_had-eta5-phi14*/	2, 124, 0, 4, 125, 0, 1, 
/* out0286_had-eta6-phi14*/	1, 124, 0, 4, 
/* out0287_had-eta7-phi14*/	0, 
/* out0288_had-eta8-phi14*/	0, 
/* out0289_had-eta9-phi14*/	5, 23, 0, 12, 23, 1, 2, 23, 2, 5, 79, 2, 3, 84, 0, 12, 
/* out0290_had-eta10-phi14*/	6, 22, 0, 4, 23, 1, 10, 23, 2, 2, 79, 2, 4, 83, 0, 11, 83, 1, 1, 
/* out0291_had-eta11-phi14*/	5, 22, 0, 8, 22, 1, 3, 22, 2, 3, 78, 2, 4, 83, 1, 9, 
/* out0292_had-eta12-phi14*/	4, 21, 0, 2, 22, 1, 8, 78, 2, 3, 82, 0, 8, 
/* out0293_had-eta13-phi14*/	4, 21, 0, 9, 21, 2, 1, 77, 2, 3, 82, 1, 7, 
/* out0294_had-eta14-phi14*/	3, 21, 1, 8, 77, 2, 4, 81, 0, 3, 
/* out0295_had-eta15-phi14*/	4, 20, 0, 5, 21, 1, 2, 81, 0, 3, 81, 1, 3, 
/* out0296_had-eta16-phi14*/	4, 20, 0, 4, 20, 1, 1, 76, 2, 3, 81, 1, 2, 
/* out0297_had-eta17-phi14*/	3, 20, 1, 5, 76, 2, 3, 80, 0, 1, 
/* out0298_had-eta18-phi14*/	3, 20, 1, 2, 76, 2, 1, 80, 0, 2, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	1, 131, 0, 2, 
/* out0301_had-eta1-phi15*/	2, 130, 0, 2, 131, 0, 6, 
/* out0302_had-eta2-phi15*/	1, 130, 0, 4, 
/* out0303_had-eta3-phi15*/	2, 129, 0, 3, 130, 0, 2, 
/* out0304_had-eta4-phi15*/	1, 129, 0, 4, 
/* out0305_had-eta5-phi15*/	2, 128, 0, 4, 129, 0, 1, 
/* out0306_had-eta6-phi15*/	1, 128, 0, 4, 
/* out0307_had-eta7-phi15*/	0, 
/* out0308_had-eta8-phi15*/	0, 
/* out0309_had-eta9-phi15*/	7, 18, 0, 1, 19, 0, 4, 19, 1, 16, 23, 0, 4, 23, 1, 1, 79, 0, 12, 79, 2, 4, 
/* out0310_had-eta10-phi15*/	6, 18, 0, 2, 18, 2, 12, 23, 1, 3, 78, 0, 1, 79, 1, 11, 79, 2, 5, 
/* out0311_had-eta11-phi15*/	8, 17, 0, 1, 17, 2, 1, 18, 1, 2, 18, 2, 4, 22, 0, 4, 22, 1, 2, 78, 0, 9, 78, 2, 5, 
/* out0312_had-eta12-phi15*/	4, 17, 2, 9, 22, 1, 2, 78, 1, 8, 78, 2, 4, 
/* out0313_had-eta13-phi15*/	5, 17, 1, 1, 17, 2, 4, 21, 0, 4, 77, 0, 7, 77, 2, 3, 
/* out0314_had-eta14-phi15*/	4, 16, 2, 4, 21, 1, 3, 77, 1, 4, 77, 2, 5, 
/* out0315_had-eta15-phi15*/	6, 16, 2, 6, 20, 0, 1, 76, 0, 3, 76, 2, 1, 77, 1, 3, 77, 2, 1, 
/* out0316_had-eta16-phi15*/	5, 16, 2, 1, 20, 0, 3, 20, 1, 1, 76, 0, 2, 76, 2, 4, 
/* out0317_had-eta17-phi15*/	4, 15, 1, 4, 20, 1, 3, 76, 1, 1, 76, 2, 3, 
/* out0318_had-eta18-phi15*/	3, 15, 1, 3, 76, 1, 2, 76, 2, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	1, 131, 0, 2, 
/* out0321_had-eta1-phi16*/	2, 130, 0, 2, 131, 0, 6, 
/* out0322_had-eta2-phi16*/	1, 130, 0, 4, 
/* out0323_had-eta3-phi16*/	2, 129, 0, 3, 130, 0, 2, 
/* out0324_had-eta4-phi16*/	1, 129, 0, 4, 
/* out0325_had-eta5-phi16*/	2, 128, 0, 4, 129, 0, 1, 
/* out0326_had-eta6-phi16*/	1, 128, 0, 4, 
/* out0327_had-eta7-phi16*/	0, 
/* out0328_had-eta8-phi16*/	1, 19, 0, 1, 
/* out0329_had-eta9-phi16*/	7, 14, 2, 7, 18, 0, 3, 19, 0, 11, 74, 0, 1, 75, 0, 5, 75, 1, 16, 79, 0, 4, 
/* out0330_had-eta10-phi16*/	6, 14, 2, 1, 18, 0, 10, 18, 1, 5, 74, 0, 2, 74, 2, 10, 79, 1, 5, 
/* out0331_had-eta11-phi16*/	8, 12, 2, 1, 17, 0, 5, 18, 1, 8, 73, 2, 1, 74, 1, 1, 74, 2, 5, 78, 0, 6, 78, 1, 2, 
/* out0332_had-eta12-phi16*/	5, 17, 0, 7, 17, 1, 3, 17, 2, 2, 73, 2, 6, 78, 1, 6, 
/* out0333_had-eta13-phi16*/	4, 16, 0, 1, 17, 1, 8, 73, 2, 2, 77, 0, 8, 
/* out0334_had-eta14-phi16*/	4, 16, 0, 7, 16, 2, 1, 77, 0, 1, 77, 1, 7, 
/* out0335_had-eta15-phi16*/	6, 16, 0, 1, 16, 1, 3, 16, 2, 3, 72, 2, 1, 76, 0, 4, 77, 1, 2, 
/* out0336_had-eta16-phi16*/	5, 15, 0, 2, 16, 1, 3, 16, 2, 1, 76, 0, 5, 76, 1, 1, 
/* out0337_had-eta17-phi16*/	3, 15, 0, 2, 15, 1, 5, 76, 1, 5, 
/* out0338_had-eta18-phi16*/	2, 15, 1, 4, 76, 1, 3, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	1, 135, 0, 2, 
/* out0341_had-eta1-phi17*/	2, 134, 0, 2, 135, 0, 6, 
/* out0342_had-eta2-phi17*/	1, 134, 0, 4, 
/* out0343_had-eta3-phi17*/	2, 133, 0, 3, 134, 0, 2, 
/* out0344_had-eta4-phi17*/	1, 133, 0, 4, 
/* out0345_had-eta5-phi17*/	2, 132, 0, 4, 133, 0, 1, 
/* out0346_had-eta6-phi17*/	1, 132, 0, 4, 
/* out0347_had-eta7-phi17*/	0, 
/* out0348_had-eta8-phi17*/	2, 14, 0, 5, 70, 0, 1, 
/* out0349_had-eta9-phi17*/	6, 14, 0, 9, 14, 1, 5, 14, 2, 6, 70, 2, 8, 74, 0, 2, 75, 0, 11, 
/* out0350_had-eta10-phi17*/	9, 12, 0, 6, 12, 2, 2, 14, 1, 6, 14, 2, 2, 18, 1, 1, 70, 2, 1, 74, 0, 11, 74, 1, 5, 74, 2, 1, 
/* out0351_had-eta11-phi17*/	5, 12, 0, 1, 12, 1, 1, 12, 2, 11, 73, 0, 5, 74, 1, 9, 
/* out0352_had-eta12-phi17*/	9, 10, 0, 1, 10, 2, 2, 12, 1, 2, 12, 2, 2, 17, 0, 3, 17, 1, 2, 73, 0, 6, 73, 1, 2, 73, 2, 4, 
/* out0353_had-eta13-phi17*/	6, 10, 2, 7, 16, 0, 1, 17, 1, 2, 72, 0, 1, 73, 1, 6, 73, 2, 3, 
/* out0354_had-eta14-phi17*/	4, 10, 2, 1, 16, 0, 6, 72, 0, 3, 72, 2, 5, 
/* out0355_had-eta15-phi17*/	2, 16, 1, 6, 72, 2, 7, 
/* out0356_had-eta16-phi17*/	7, 9, 2, 1, 15, 0, 2, 16, 1, 3, 71, 2, 1, 72, 2, 2, 76, 0, 2, 76, 1, 1, 
/* out0357_had-eta17-phi17*/	3, 15, 0, 5, 71, 2, 3, 76, 1, 2, 
/* out0358_had-eta18-phi17*/	3, 15, 0, 1, 71, 2, 3, 76, 1, 1, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	1, 135, 0, 2, 
/* out0361_had-eta1-phi18*/	2, 134, 0, 2, 135, 0, 6, 
/* out0362_had-eta2-phi18*/	1, 134, 0, 4, 
/* out0363_had-eta3-phi18*/	2, 133, 0, 3, 134, 0, 2, 
/* out0364_had-eta4-phi18*/	1, 133, 0, 4, 
/* out0365_had-eta5-phi18*/	2, 132, 0, 4, 133, 0, 1, 
/* out0366_had-eta6-phi18*/	1, 132, 0, 4, 
/* out0367_had-eta7-phi18*/	0, 
/* out0368_had-eta8-phi18*/	0, 
/* out0369_had-eta9-phi18*/	7, 13, 0, 4, 13, 2, 5, 14, 0, 2, 14, 1, 4, 70, 0, 14, 70, 1, 6, 70, 2, 5, 
/* out0370_had-eta10-phi18*/	8, 12, 0, 6, 13, 2, 9, 14, 1, 1, 68, 0, 6, 68, 2, 3, 70, 1, 5, 70, 2, 2, 74, 1, 1, 
/* out0371_had-eta11-phi18*/	5, 11, 2, 1, 12, 0, 3, 12, 1, 10, 68, 2, 12, 73, 0, 1, 
/* out0372_had-eta12-phi18*/	7, 10, 0, 8, 12, 1, 3, 67, 2, 2, 68, 1, 1, 68, 2, 1, 73, 0, 4, 73, 1, 4, 
/* out0373_had-eta13-phi18*/	6, 10, 0, 3, 10, 1, 3, 10, 2, 4, 67, 2, 3, 72, 0, 2, 73, 1, 4, 
/* out0374_had-eta14-phi18*/	5, 9, 0, 2, 10, 1, 4, 10, 2, 2, 72, 0, 8, 72, 1, 1, 
/* out0375_had-eta15-phi18*/	5, 9, 0, 1, 9, 2, 5, 16, 1, 1, 72, 1, 6, 72, 2, 1, 
/* out0376_had-eta16-phi18*/	3, 9, 2, 5, 71, 0, 3, 72, 1, 3, 
/* out0377_had-eta17-phi18*/	4, 9, 2, 1, 15, 0, 4, 71, 0, 2, 71, 2, 4, 
/* out0378_had-eta18-phi18*/	1, 71, 2, 5, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	1, 139, 0, 2, 
/* out0381_had-eta1-phi19*/	2, 138, 0, 2, 139, 0, 6, 
/* out0382_had-eta2-phi19*/	1, 138, 0, 4, 
/* out0383_had-eta3-phi19*/	2, 137, 0, 3, 138, 0, 2, 
/* out0384_had-eta4-phi19*/	1, 137, 0, 4, 
/* out0385_had-eta5-phi19*/	2, 136, 0, 4, 137, 0, 1, 
/* out0386_had-eta6-phi19*/	1, 136, 0, 4, 
/* out0387_had-eta7-phi19*/	0, 
/* out0388_had-eta8-phi19*/	0, 
/* out0389_had-eta9-phi19*/	6, 13, 0, 12, 13, 1, 3, 69, 0, 5, 69, 2, 8, 70, 0, 1, 70, 1, 4, 
/* out0390_had-eta10-phi19*/	7, 11, 0, 3, 13, 1, 12, 13, 2, 2, 68, 0, 9, 68, 1, 1, 69, 2, 7, 70, 1, 1, 
/* out0391_had-eta11-phi19*/	4, 11, 0, 5, 11, 2, 8, 68, 0, 1, 68, 1, 13, 
/* out0392_had-eta12-phi19*/	6, 10, 0, 3, 11, 1, 2, 11, 2, 7, 67, 0, 9, 67, 2, 2, 68, 1, 1, 
/* out0393_had-eta13-phi19*/	6, 10, 0, 1, 10, 1, 6, 48, 2, 2, 67, 0, 1, 67, 1, 2, 67, 2, 7, 
/* out0394_had-eta14-phi19*/	8, 9, 0, 4, 10, 1, 3, 48, 2, 1, 61, 2, 1, 67, 1, 1, 67, 2, 2, 72, 0, 2, 72, 1, 2, 
/* out0395_had-eta15-phi19*/	5, 9, 0, 5, 9, 1, 1, 9, 2, 1, 61, 2, 3, 72, 1, 4, 
/* out0396_had-eta16-phi19*/	4, 9, 1, 3, 9, 2, 2, 61, 2, 1, 71, 0, 4, 
/* out0397_had-eta17-phi19*/	4, 9, 1, 2, 9, 2, 1, 71, 0, 4, 71, 1, 1, 
/* out0398_had-eta18-phi19*/	1, 71, 1, 5, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	1, 139, 0, 2, 
/* out0401_had-eta1-phi20*/	2, 138, 0, 2, 139, 0, 6, 
/* out0402_had-eta2-phi20*/	1, 138, 0, 4, 
/* out0403_had-eta3-phi20*/	2, 137, 0, 3, 138, 0, 2, 
/* out0404_had-eta4-phi20*/	1, 137, 0, 4, 
/* out0405_had-eta5-phi20*/	2, 136, 0, 4, 137, 0, 1, 
/* out0406_had-eta6-phi20*/	1, 136, 0, 4, 
/* out0407_had-eta7-phi20*/	0, 
/* out0408_had-eta8-phi20*/	0, 
/* out0409_had-eta9-phi20*/	5, 13, 1, 1, 51, 0, 8, 51, 2, 3, 69, 0, 11, 69, 1, 7, 
/* out0410_had-eta10-phi20*/	6, 11, 0, 2, 51, 2, 13, 65, 0, 6, 65, 2, 1, 69, 1, 9, 69, 2, 1, 
/* out0411_had-eta11-phi20*/	4, 11, 0, 6, 11, 1, 7, 65, 0, 2, 65, 2, 12, 
/* out0412_had-eta12-phi20*/	5, 11, 1, 7, 48, 0, 4, 65, 2, 3, 67, 0, 6, 67, 1, 2, 
/* out0413_had-eta13-phi20*/	3, 48, 0, 4, 48, 2, 6, 67, 1, 10, 
/* out0414_had-eta14-phi20*/	4, 9, 0, 1, 48, 2, 7, 61, 0, 6, 67, 1, 1, 
/* out0415_had-eta15-phi20*/	4, 9, 0, 3, 9, 1, 4, 61, 0, 1, 61, 2, 6, 
/* out0416_had-eta16-phi20*/	3, 9, 1, 5, 61, 2, 5, 71, 0, 1, 
/* out0417_had-eta17-phi20*/	3, 9, 1, 1, 71, 0, 2, 71, 1, 4, 
/* out0418_had-eta18-phi20*/	1, 71, 1, 5, 
/* out0419_had-eta19-phi20*/	1, 71, 1, 1, 
/* out0420_had-eta0-phi21*/	1, 143, 0, 2, 
/* out0421_had-eta1-phi21*/	2, 142, 0, 2, 143, 0, 6, 
/* out0422_had-eta2-phi21*/	1, 142, 0, 4, 
/* out0423_had-eta3-phi21*/	2, 141, 0, 3, 142, 0, 2, 
/* out0424_had-eta4-phi21*/	1, 141, 0, 4, 
/* out0425_had-eta5-phi21*/	2, 140, 0, 4, 141, 0, 1, 
/* out0426_had-eta6-phi21*/	1, 140, 0, 4, 
/* out0427_had-eta7-phi21*/	0, 
/* out0428_had-eta8-phi21*/	0, 
/* out0429_had-eta9-phi21*/	5, 50, 2, 1, 51, 0, 8, 51, 1, 3, 66, 0, 11, 66, 2, 7, 
/* out0430_had-eta10-phi21*/	6, 49, 0, 2, 51, 1, 13, 65, 0, 6, 65, 1, 1, 66, 1, 1, 66, 2, 9, 
/* out0431_had-eta11-phi21*/	4, 49, 0, 6, 49, 2, 7, 65, 0, 2, 65, 1, 12, 
/* out0432_had-eta12-phi21*/	5, 48, 0, 4, 49, 2, 7, 62, 0, 6, 62, 2, 2, 65, 1, 3, 
/* out0433_had-eta13-phi21*/	3, 48, 0, 4, 48, 1, 6, 62, 2, 10, 
/* out0434_had-eta14-phi21*/	4, 5, 0, 1, 48, 1, 7, 61, 0, 7, 62, 2, 1, 
/* out0435_had-eta15-phi21*/	4, 5, 0, 3, 5, 2, 4, 61, 0, 1, 61, 1, 6, 
/* out0436_had-eta16-phi21*/	3, 5, 2, 5, 56, 0, 1, 61, 1, 5, 
/* out0437_had-eta17-phi21*/	3, 5, 2, 1, 56, 0, 2, 56, 2, 4, 
/* out0438_had-eta18-phi21*/	1, 56, 2, 5, 
/* out0439_had-eta19-phi21*/	1, 56, 2, 1, 
/* out0440_had-eta0-phi22*/	1, 143, 0, 2, 
/* out0441_had-eta1-phi22*/	2, 142, 0, 2, 143, 0, 6, 
/* out0442_had-eta2-phi22*/	1, 142, 0, 4, 
/* out0443_had-eta3-phi22*/	2, 141, 0, 3, 142, 0, 2, 
/* out0444_had-eta4-phi22*/	1, 141, 0, 4, 
/* out0445_had-eta5-phi22*/	2, 140, 0, 4, 141, 0, 1, 
/* out0446_had-eta6-phi22*/	1, 140, 0, 4, 
/* out0447_had-eta7-phi22*/	0, 
/* out0448_had-eta8-phi22*/	0, 
/* out0449_had-eta9-phi22*/	6, 50, 0, 12, 50, 2, 3, 64, 0, 1, 64, 2, 4, 66, 0, 5, 66, 1, 8, 
/* out0450_had-eta10-phi22*/	7, 49, 0, 3, 50, 1, 2, 50, 2, 12, 63, 0, 9, 63, 2, 1, 64, 2, 1, 66, 1, 7, 
/* out0451_had-eta11-phi22*/	4, 49, 0, 5, 49, 1, 8, 63, 0, 1, 63, 2, 13, 
/* out0452_had-eta12-phi22*/	6, 6, 0, 3, 49, 1, 7, 49, 2, 2, 62, 0, 9, 62, 1, 2, 63, 2, 1, 
/* out0453_had-eta13-phi22*/	6, 6, 0, 1, 6, 2, 6, 48, 1, 2, 62, 0, 1, 62, 1, 7, 62, 2, 2, 
/* out0454_had-eta14-phi22*/	9, 5, 0, 4, 6, 2, 3, 48, 1, 1, 57, 0, 2, 57, 2, 2, 61, 0, 1, 61, 1, 1, 62, 1, 2, 62, 2, 1, 
/* out0455_had-eta15-phi22*/	5, 5, 0, 5, 5, 1, 1, 5, 2, 1, 57, 2, 4, 61, 1, 3, 
/* out0456_had-eta16-phi22*/	4, 5, 1, 2, 5, 2, 3, 56, 0, 4, 61, 1, 1, 
/* out0457_had-eta17-phi22*/	4, 5, 1, 1, 5, 2, 2, 56, 0, 4, 56, 2, 1, 
/* out0458_had-eta18-phi22*/	1, 56, 2, 5, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	1, 147, 0, 2, 
/* out0461_had-eta1-phi23*/	2, 146, 0, 2, 147, 0, 6, 
/* out0462_had-eta2-phi23*/	1, 146, 0, 4, 
/* out0463_had-eta3-phi23*/	2, 145, 0, 3, 146, 0, 2, 
/* out0464_had-eta4-phi23*/	1, 145, 0, 4, 
/* out0465_had-eta5-phi23*/	2, 144, 0, 4, 145, 0, 1, 
/* out0466_had-eta6-phi23*/	1, 144, 0, 4, 
/* out0467_had-eta7-phi23*/	0, 
/* out0468_had-eta8-phi23*/	0, 
/* out0469_had-eta9-phi23*/	7, 8, 0, 2, 8, 2, 4, 50, 0, 4, 50, 1, 5, 64, 0, 14, 64, 1, 5, 64, 2, 6, 
/* out0470_had-eta10-phi23*/	8, 7, 0, 6, 8, 2, 1, 50, 1, 9, 59, 2, 1, 63, 0, 6, 63, 1, 3, 64, 1, 2, 64, 2, 5, 
/* out0471_had-eta11-phi23*/	5, 7, 0, 3, 7, 2, 10, 49, 1, 1, 58, 0, 1, 63, 1, 12, 
/* out0472_had-eta12-phi23*/	7, 6, 0, 8, 7, 2, 3, 58, 0, 4, 58, 2, 4, 62, 1, 2, 63, 1, 1, 63, 2, 1, 
/* out0473_had-eta13-phi23*/	6, 6, 0, 3, 6, 1, 4, 6, 2, 3, 57, 0, 2, 58, 2, 4, 62, 1, 3, 
/* out0474_had-eta14-phi23*/	5, 5, 0, 2, 6, 1, 2, 6, 2, 4, 57, 0, 8, 57, 2, 1, 
/* out0475_had-eta15-phi23*/	5, 1, 2, 1, 5, 0, 1, 5, 1, 5, 57, 1, 1, 57, 2, 6, 
/* out0476_had-eta16-phi23*/	3, 5, 1, 5, 56, 0, 3, 57, 2, 3, 
/* out0477_had-eta17-phi23*/	4, 0, 0, 4, 5, 1, 1, 56, 0, 2, 56, 1, 4, 
/* out0478_had-eta18-phi23*/	1, 56, 1, 5, 
/* out0479_had-eta19-phi23*/	0, 
/* out0480_had-eta0-phi24*/	1, 147, 0, 2, 
/* out0481_had-eta1-phi24*/	2, 146, 0, 2, 147, 0, 6, 
/* out0482_had-eta2-phi24*/	1, 146, 0, 4, 
/* out0483_had-eta3-phi24*/	2, 145, 0, 3, 146, 0, 2, 
/* out0484_had-eta4-phi24*/	1, 145, 0, 4, 
/* out0485_had-eta5-phi24*/	2, 144, 0, 4, 145, 0, 1, 
/* out0486_had-eta6-phi24*/	1, 144, 0, 4, 
/* out0487_had-eta7-phi24*/	0, 
/* out0488_had-eta8-phi24*/	2, 8, 0, 5, 64, 0, 1, 
/* out0489_had-eta9-phi24*/	6, 8, 0, 9, 8, 1, 6, 8, 2, 5, 59, 0, 2, 60, 1, 11, 64, 1, 8, 
/* out0490_had-eta10-phi24*/	9, 3, 2, 1, 7, 0, 6, 7, 1, 2, 8, 1, 2, 8, 2, 6, 59, 0, 11, 59, 1, 1, 59, 2, 5, 64, 1, 1, 
/* out0491_had-eta11-phi24*/	5, 7, 0, 1, 7, 1, 11, 7, 2, 1, 58, 0, 5, 59, 2, 9, 
/* out0492_had-eta12-phi24*/	9, 2, 0, 3, 2, 2, 2, 6, 0, 1, 6, 1, 2, 7, 1, 2, 7, 2, 2, 58, 0, 6, 58, 1, 4, 58, 2, 2, 
/* out0493_had-eta13-phi24*/	6, 1, 0, 1, 2, 2, 2, 6, 1, 7, 57, 0, 1, 58, 1, 3, 58, 2, 6, 
/* out0494_had-eta14-phi24*/	4, 1, 0, 6, 6, 1, 1, 57, 0, 3, 57, 1, 5, 
/* out0495_had-eta15-phi24*/	2, 1, 2, 6, 57, 1, 7, 
/* out0496_had-eta16-phi24*/	7, 0, 0, 2, 1, 2, 3, 5, 1, 1, 52, 0, 2, 52, 2, 1, 56, 1, 1, 57, 1, 2, 
/* out0497_had-eta17-phi24*/	3, 0, 0, 5, 52, 2, 2, 56, 1, 3, 
/* out0498_had-eta18-phi24*/	3, 0, 0, 1, 52, 2, 1, 56, 1, 3, 
/* out0499_had-eta19-phi24*/	0, 
/* out0500_had-eta0-phi25*/	1, 151, 0, 2, 
/* out0501_had-eta1-phi25*/	2, 150, 0, 2, 151, 0, 6, 
/* out0502_had-eta2-phi25*/	1, 150, 0, 4, 
/* out0503_had-eta3-phi25*/	2, 149, 0, 3, 150, 0, 2, 
/* out0504_had-eta4-phi25*/	1, 149, 0, 4, 
/* out0505_had-eta5-phi25*/	2, 148, 0, 4, 149, 0, 1, 
/* out0506_had-eta6-phi25*/	1, 148, 0, 4, 
/* out0507_had-eta7-phi25*/	0, 
/* out0508_had-eta8-phi25*/	1, 4, 1, 1, 
/* out0509_had-eta9-phi25*/	7, 3, 0, 3, 4, 1, 11, 8, 1, 7, 55, 0, 4, 59, 0, 1, 60, 0, 16, 60, 1, 5, 
/* out0510_had-eta10-phi25*/	6, 3, 0, 10, 3, 2, 5, 8, 1, 1, 55, 2, 5, 59, 0, 2, 59, 1, 10, 
/* out0511_had-eta11-phi25*/	8, 2, 0, 5, 3, 2, 8, 7, 1, 1, 54, 0, 6, 54, 2, 2, 58, 1, 1, 59, 1, 5, 59, 2, 1, 
/* out0512_had-eta12-phi25*/	5, 2, 0, 7, 2, 1, 2, 2, 2, 3, 54, 2, 6, 58, 1, 6, 
/* out0513_had-eta13-phi25*/	4, 1, 0, 1, 2, 2, 8, 53, 0, 8, 58, 1, 2, 
/* out0514_had-eta14-phi25*/	4, 1, 0, 7, 1, 1, 1, 53, 0, 1, 53, 2, 7, 
/* out0515_had-eta15-phi25*/	6, 1, 0, 1, 1, 1, 3, 1, 2, 3, 52, 0, 4, 53, 2, 2, 57, 1, 1, 
/* out0516_had-eta16-phi25*/	5, 0, 0, 2, 1, 1, 1, 1, 2, 3, 52, 0, 5, 52, 2, 1, 
/* out0517_had-eta17-phi25*/	3, 0, 0, 2, 0, 1, 5, 52, 2, 5, 
/* out0518_had-eta18-phi25*/	2, 0, 1, 4, 52, 2, 3, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	1, 151, 0, 2, 
/* out0521_had-eta1-phi26*/	2, 150, 0, 2, 151, 0, 6, 
/* out0522_had-eta2-phi26*/	1, 150, 0, 4, 
/* out0523_had-eta3-phi26*/	2, 149, 0, 3, 150, 0, 2, 
/* out0524_had-eta4-phi26*/	1, 149, 0, 4, 
/* out0525_had-eta5-phi26*/	2, 148, 0, 4, 149, 0, 1, 
/* out0526_had-eta6-phi26*/	1, 148, 0, 4, 
/* out0527_had-eta7-phi26*/	0, 
/* out0528_had-eta8-phi26*/	0, 
/* out0529_had-eta9-phi26*/	5, 3, 0, 1, 4, 0, 16, 4, 1, 4, 55, 0, 12, 55, 1, 4, 
/* out0530_had-eta10-phi26*/	5, 3, 0, 2, 3, 1, 12, 54, 0, 1, 55, 1, 5, 55, 2, 11, 
/* out0531_had-eta11-phi26*/	6, 2, 0, 1, 2, 1, 1, 3, 1, 4, 3, 2, 2, 54, 0, 9, 54, 1, 5, 
/* out0532_had-eta12-phi26*/	3, 2, 1, 9, 54, 1, 4, 54, 2, 8, 
/* out0533_had-eta13-phi26*/	4, 2, 1, 4, 2, 2, 1, 53, 0, 7, 53, 1, 3, 
/* out0534_had-eta14-phi26*/	3, 1, 1, 4, 53, 1, 5, 53, 2, 4, 
/* out0535_had-eta15-phi26*/	5, 1, 1, 6, 52, 0, 3, 52, 1, 1, 53, 1, 1, 53, 2, 3, 
/* out0536_had-eta16-phi26*/	3, 1, 1, 1, 52, 0, 2, 52, 1, 4, 
/* out0537_had-eta17-phi26*/	3, 0, 1, 4, 52, 1, 3, 52, 2, 1, 
/* out0538_had-eta18-phi26*/	3, 0, 1, 3, 52, 1, 1, 52, 2, 2, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	1, 55, 1, 3, 
/* out0550_had-eta10-phi27*/	1, 55, 1, 4, 
/* out0551_had-eta11-phi27*/	1, 54, 1, 4, 
/* out0552_had-eta12-phi27*/	1, 54, 1, 3, 
/* out0553_had-eta13-phi27*/	1, 53, 1, 3, 
/* out0554_had-eta14-phi27*/	1, 53, 1, 4, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	1, 52, 1, 3, 
/* out0557_had-eta17-phi27*/	1, 52, 1, 3, 
/* out0558_had-eta18-phi27*/	1, 52, 1, 1, 
/* out0559_had-eta19-phi27*/	0, 
};