parameter integer matrixH [0:7121] = {
/* num inputs = 140(in0-in139) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2213 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	4,79,0,16,79,1,11,79,2,3,89,2,3,
/* out0006_em-eta6-phi0*/	6,68,0,10,68,1,4,79,1,4,79,2,13,80,0,1,80,2,1,
/* out0007_em-eta7-phi0*/	4,57,0,5,68,0,6,68,1,8,68,2,16,
/* out0008_em-eta8-phi0*/	4,57,0,11,57,1,6,57,2,3,273,2,3,
/* out0009_em-eta9-phi0*/	7,46,0,6,57,1,2,57,2,10,265,0,1,265,1,2,273,1,4,273,2,10,
/* out0010_em-eta10-phi0*/	5,46,0,7,46,1,3,46,2,7,265,0,12,265,1,1,
/* out0011_em-eta11-phi0*/	7,35,0,4,46,2,8,131,2,5,257,0,1,257,1,2,265,0,3,265,2,2,
/* out0012_em-eta12-phi0*/	8,35,0,8,35,1,1,35,2,1,124,0,1,124,1,1,131,1,2,131,2,7,257,0,9,
/* out0013_em-eta13-phi0*/	5,35,2,8,124,0,9,249,1,1,257,0,4,257,2,1,
/* out0014_em-eta14-phi0*/	5,24,0,8,35,2,4,124,0,5,124,2,1,249,0,5,
/* out0015_em-eta15-phi0*/	4,24,0,4,24,2,2,117,0,4,249,0,5,
/* out0016_em-eta16-phi0*/	3,24,2,5,117,0,5,249,0,1,
/* out0017_em-eta17-phi0*/	4,14,2,3,24,2,2,117,0,2,242,2,3,
/* out0018_em-eta18-phi0*/	4,14,2,5,111,2,2,242,0,1,242,2,1,
/* out0019_em-eta19-phi0*/	4,14,0,2,14,2,1,111,0,1,111,2,2,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	6,79,1,1,80,0,7,80,1,1,89,1,14,89,2,13,90,0,1,
/* out0026_em-eta6-phi1*/	4,68,1,1,80,0,8,80,1,5,80,2,14,
/* out0027_em-eta7-phi1*/	5,68,1,3,69,0,15,69,1,1,69,2,3,80,2,1,
/* out0028_em-eta8-phi1*/	6,57,1,6,58,0,4,69,2,10,273,1,1,273,2,2,274,0,1,
/* out0029_em-eta9-phi1*/	10,46,0,3,46,1,1,57,1,2,57,2,3,58,0,7,58,2,5,265,1,4,273,1,11,273,2,1,274,0,7,
/* out0030_em-eta10-phi1*/	5,46,1,9,47,0,2,58,2,3,265,1,9,265,2,7,
/* out0031_em-eta11-phi1*/	11,35,0,1,35,1,1,46,1,3,46,2,1,47,0,4,47,2,2,131,1,2,131,2,4,257,1,6,265,2,6,266,0,1,
/* out0032_em-eta12-phi1*/	9,35,0,3,35,1,8,47,2,1,124,1,4,131,1,11,132,0,1,257,0,2,257,1,6,257,2,3,
/* out0033_em-eta13-phi1*/	8,35,1,5,35,2,2,36,0,1,124,0,1,124,1,8,124,2,2,249,1,2,257,2,7,
/* out0034_em-eta14-phi1*/	8,24,0,3,24,1,3,35,2,1,36,2,1,117,1,1,124,2,8,249,0,2,249,1,6,
/* out0035_em-eta15-phi1*/	7,24,0,1,24,1,5,24,2,1,117,0,1,117,1,7,249,0,3,249,2,3,
/* out0036_em-eta16-phi1*/	7,24,1,2,24,2,3,117,0,3,117,1,1,117,2,3,242,2,3,249,2,3,
/* out0037_em-eta17-phi1*/	6,14,2,3,24,2,2,111,2,1,117,0,1,117,2,4,242,2,6,
/* out0038_em-eta18-phi1*/	4,14,0,3,14,2,2,111,2,6,242,0,2,
/* out0039_em-eta19-phi1*/	3,14,0,2,111,0,2,111,2,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	5,80,1,1,89,1,2,90,0,15,90,1,10,90,2,11,
/* out0046_em-eta6-phi2*/	4,80,1,9,81,0,14,81,2,2,90,2,4,
/* out0047_em-eta7-phi2*/	4,69,0,1,69,1,12,70,0,2,81,2,8,
/* out0048_em-eta8-phi2*/	9,58,0,3,58,1,3,69,1,3,69,2,3,70,0,4,70,2,3,274,1,7,280,0,1,280,1,1,
/* out0049_em-eta9-phi2*/	6,58,0,2,58,1,10,58,2,4,274,0,7,274,1,6,274,2,6,
/* out0050_em-eta10-phi2*/	9,47,0,7,47,1,2,58,1,1,58,2,4,265,2,1,266,0,3,266,1,6,274,0,1,274,2,4,
/* out0051_em-eta11-phi2*/	9,47,0,3,47,1,2,47,2,5,131,1,1,132,0,2,132,1,6,266,0,11,266,1,1,266,2,2,
/* out0052_em-eta12-phi2*/	12,35,1,1,36,0,3,47,2,6,132,0,11,132,1,1,132,2,1,257,1,2,257,2,3,258,0,2,258,1,1,266,0,1,266,2,1,
/* out0053_em-eta13-phi2*/	10,36,0,7,124,1,3,124,2,2,125,0,1,125,1,1,132,0,2,132,2,2,249,1,1,257,2,2,258,0,7,
/* out0054_em-eta14-phi2*/	7,24,1,1,36,2,6,124,2,3,125,0,7,249,1,6,249,2,1,258,0,1,
/* out0055_em-eta15-phi2*/	6,24,1,3,25,0,1,36,2,1,117,1,6,125,0,2,249,2,6,
/* out0056_em-eta16-phi2*/	8,24,1,2,25,0,3,117,1,1,117,2,6,242,0,1,242,2,2,249,2,2,250,0,1,
/* out0057_em-eta17-phi2*/	11,14,0,2,14,2,2,24,2,1,25,0,1,25,2,2,111,0,1,111,2,2,117,2,3,118,0,1,242,0,5,242,2,1,
/* out0058_em-eta18-phi2*/	4,14,0,4,111,0,5,111,2,2,242,0,1,
/* out0059_em-eta19-phi2*/	2,14,0,1,111,0,2,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	0,
/* out0065_em-eta5-phi3*/	3,90,1,6,91,0,15,91,2,2,
/* out0066_em-eta6-phi3*/	6,81,0,2,81,1,14,81,2,1,82,0,3,90,2,1,91,2,8,
/* out0067_em-eta7-phi3*/	6,70,0,7,70,1,5,81,1,2,81,2,5,82,0,2,82,2,2,
/* out0068_em-eta8-phi3*/	7,70,0,3,70,1,5,70,2,11,274,1,1,280,0,12,280,1,7,280,2,9,
/* out0069_em-eta9-phi3*/	10,58,1,2,59,0,13,70,2,2,274,1,2,274,2,5,275,0,6,275,1,4,280,0,2,280,1,7,280,2,5,
/* out0070_em-eta10-phi3*/	6,47,1,3,59,0,1,59,2,9,266,1,8,274,2,1,275,0,7,
/* out0071_em-eta11-phi3*/	9,47,1,8,48,0,3,132,1,6,137,0,10,137,1,7,137,2,3,266,1,1,266,2,11,267,0,1,
/* out0072_em-eta12-phi3*/	11,36,0,3,36,1,2,47,1,1,47,2,2,48,0,1,48,2,1,132,1,3,132,2,10,133,0,1,258,1,9,266,2,2,
/* out0073_em-eta13-phi3*/	7,36,0,2,36,1,5,125,1,8,132,2,3,258,0,4,258,1,2,258,2,4,
/* out0074_em-eta14-phi3*/	8,36,1,1,36,2,6,125,0,4,125,1,3,125,2,3,250,1,2,258,0,2,258,2,3,
/* out0075_em-eta15-phi3*/	8,25,0,4,36,2,1,118,1,1,125,0,2,125,2,4,249,2,1,250,0,5,250,1,1,
/* out0076_em-eta16-phi3*/	5,25,0,4,118,0,5,118,1,1,242,0,1,250,0,5,
/* out0077_em-eta17-phi3*/	4,25,2,4,118,0,5,242,0,5,250,0,1,
/* out0078_em-eta18-phi3*/	4,14,0,2,25,2,2,111,0,4,118,0,1,
/* out0079_em-eta19-phi3*/	1,111,0,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	0,
/* out0085_em-eta5-phi4*/	7,91,0,1,91,1,14,91,2,1,92,0,6,97,0,15,97,1,14,97,2,12,
/* out0086_em-eta6-phi4*/	6,82,0,9,82,1,7,91,1,2,91,2,5,92,0,2,92,2,3,
/* out0087_em-eta7-phi4*/	5,70,1,1,71,0,3,82,0,2,82,1,3,82,2,14,
/* out0088_em-eta8-phi4*/	8,70,1,5,71,0,10,71,2,4,280,0,1,280,1,1,280,2,2,281,0,2,281,2,1,
/* out0089_em-eta9-phi4*/	9,59,0,2,59,1,12,71,2,2,275,0,1,275,1,12,275,2,4,281,0,6,281,1,5,281,2,1,
/* out0090_em-eta10-phi4*/	6,48,0,2,59,1,4,59,2,7,267,1,4,275,0,2,275,2,10,
/* out0091_em-eta11-phi4*/	9,48,0,10,48,1,1,48,2,1,133,1,2,137,0,6,137,1,9,137,2,13,267,0,9,267,1,4,
/* out0092_em-eta12-phi4*/	7,36,1,1,48,2,8,133,0,8,133,1,6,258,1,4,267,0,6,267,2,1,
/* out0093_em-eta13-phi4*/	8,36,1,5,37,0,2,48,2,1,125,1,3,133,0,7,133,2,1,258,2,7,259,0,2,
/* out0094_em-eta14-phi4*/	10,36,1,2,36,2,1,37,0,2,37,2,1,125,1,1,125,2,6,126,0,2,250,1,5,258,2,2,259,0,1,
/* out0095_em-eta15-phi4*/	8,25,0,2,25,1,3,118,1,4,125,2,3,126,0,1,250,0,1,250,1,4,250,2,1,
/* out0096_em-eta16-phi4*/	7,25,0,1,25,1,3,118,0,1,118,1,6,118,2,1,250,0,2,250,2,3,
/* out0097_em-eta17-phi4*/	5,25,2,4,118,0,2,118,2,3,250,0,1,250,2,2,
/* out0098_em-eta18-phi4*/	3,25,2,2,118,0,1,118,2,2,
/* out0099_em-eta19-phi4*/	0,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	0,
/* out0105_em-eta5-phi5*/	8,92,0,8,92,1,13,97,0,1,97,1,2,97,2,4,98,0,12,98,1,8,98,2,4,
/* out0106_em-eta6-phi5*/	4,82,1,3,83,0,9,92,1,3,92,2,13,
/* out0107_em-eta7-phi5*/	5,71,0,1,71,1,3,82,1,3,83,0,7,83,2,8,
/* out0108_em-eta8-phi5*/	3,71,0,2,71,1,13,71,2,5,
/* out0109_em-eta9-phi5*/	8,60,0,11,71,2,5,275,2,1,276,0,4,276,1,8,281,0,8,281,1,11,281,2,14,
/* out0110_em-eta10-phi5*/	6,48,1,1,60,0,5,60,2,7,267,1,3,275,2,1,276,0,12,
/* out0111_em-eta11-phi5*/	8,48,1,11,60,2,1,133,1,2,138,0,10,138,1,6,138,2,4,267,1,5,267,2,9,
/* out0112_em-eta12-phi5*/	9,37,0,1,48,1,3,48,2,5,133,1,6,133,2,7,138,0,2,138,1,2,259,1,5,267,2,6,
/* out0113_em-eta13-phi5*/	5,37,0,8,126,1,4,133,2,8,259,0,7,259,1,3,
/* out0114_em-eta14-phi5*/	6,37,0,3,37,2,4,126,0,5,126,1,4,250,1,2,259,0,6,
/* out0115_em-eta15-phi5*/	6,25,1,3,37,2,3,118,1,1,126,0,7,250,1,2,250,2,4,
/* out0116_em-eta16-phi5*/	5,25,1,5,118,1,3,118,2,3,126,0,1,250,2,5,
/* out0117_em-eta17-phi5*/	4,25,1,2,25,2,1,118,2,6,250,2,1,
/* out0118_em-eta18-phi5*/	2,25,2,1,118,2,1,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	0,
/* out0125_em-eta5-phi6*/	8,93,0,13,93,1,8,98,0,4,98,1,8,98,2,12,99,0,4,99,1,2,99,2,1,
/* out0126_em-eta6-phi6*/	4,83,1,9,84,0,3,93,0,3,93,2,13,
/* out0127_em-eta7-phi6*/	5,72,0,3,72,1,1,83,1,7,83,2,8,84,0,3,
/* out0128_em-eta8-phi6*/	3,72,0,13,72,1,2,72,2,5,
/* out0129_em-eta9-phi6*/	8,60,1,11,72,2,5,276,1,8,276,2,4,277,0,1,282,0,14,282,1,11,282,2,8,
/* out0130_em-eta10-phi6*/	6,49,0,1,60,1,5,60,2,7,268,1,3,276,2,12,277,0,1,
/* out0131_em-eta11-phi6*/	8,49,0,11,60,2,1,134,1,2,138,0,4,138,1,6,138,2,10,268,0,9,268,1,5,
/* out0132_em-eta12-phi6*/	9,37,1,1,49,0,3,49,2,5,134,0,7,134,1,6,138,1,2,138,2,2,259,1,5,268,0,6,
/* out0133_em-eta13-phi6*/	5,37,1,8,126,1,4,134,0,8,259,1,3,259,2,7,
/* out0134_em-eta14-phi6*/	6,37,1,3,37,2,4,126,1,4,126,2,5,251,1,2,259,2,6,
/* out0135_em-eta15-phi6*/	6,26,0,3,37,2,3,119,1,1,126,2,7,251,0,4,251,1,2,
/* out0136_em-eta16-phi6*/	5,26,0,5,119,0,3,119,1,3,126,2,1,251,0,5,
/* out0137_em-eta17-phi6*/	4,26,0,2,26,2,1,119,0,6,251,0,1,
/* out0138_em-eta18-phi6*/	2,26,2,1,119,0,1,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	0,
/* out0145_em-eta5-phi7*/	7,93,1,6,94,0,14,94,1,1,94,2,1,99,0,12,99,1,14,99,2,15,
/* out0146_em-eta6-phi7*/	6,84,0,7,84,1,9,93,1,2,93,2,3,94,0,2,94,2,5,
/* out0147_em-eta7-phi7*/	5,72,1,3,73,0,1,84,0,3,84,1,2,84,2,14,
/* out0148_em-eta8-phi7*/	8,72,1,10,72,2,4,73,0,5,282,0,1,282,2,2,283,0,2,283,1,1,283,2,1,
/* out0149_em-eta9-phi7*/	9,61,0,12,61,1,2,72,2,2,277,0,4,277,1,12,277,2,1,282,0,1,282,1,5,282,2,6,
/* out0150_em-eta10-phi7*/	6,49,1,2,61,0,4,61,2,7,268,1,4,277,0,10,277,2,1,
/* out0151_em-eta11-phi7*/	9,49,0,1,49,1,10,49,2,1,134,1,2,139,0,13,139,1,9,139,2,6,268,1,4,268,2,9,
/* out0152_em-eta12-phi7*/	7,38,0,1,49,2,8,134,1,6,134,2,8,260,1,4,268,0,1,268,2,6,
/* out0153_em-eta13-phi7*/	8,37,1,2,38,0,5,49,2,1,127,1,3,134,0,1,134,2,7,259,2,2,260,0,7,
/* out0154_em-eta14-phi7*/	10,37,1,2,37,2,1,38,0,2,38,2,1,126,2,2,127,0,6,127,1,1,251,1,5,259,2,1,260,0,2,
/* out0155_em-eta15-phi7*/	8,26,0,3,26,1,2,119,1,4,126,2,1,127,0,3,251,0,1,251,1,4,251,2,1,
/* out0156_em-eta16-phi7*/	7,26,0,3,26,1,1,119,0,1,119,1,6,119,2,1,251,0,3,251,2,2,
/* out0157_em-eta17-phi7*/	5,26,2,4,119,0,3,119,2,2,251,0,2,251,2,1,
/* out0158_em-eta18-phi7*/	3,26,2,2,119,0,2,119,2,1,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	0,
/* out0165_em-eta5-phi8*/	5,94,1,15,94,2,2,95,0,13,95,1,2,95,2,1,
/* out0166_em-eta6-phi8*/	5,84,1,3,85,0,14,85,1,2,85,2,1,94,2,8,
/* out0167_em-eta7-phi8*/	6,73,0,5,73,1,7,84,1,2,84,2,2,85,0,2,85,2,5,
/* out0168_em-eta8-phi8*/	7,73,0,5,73,1,3,73,2,11,278,1,1,283,0,9,283,1,7,283,2,12,
/* out0169_em-eta9-phi8*/	10,61,1,13,62,0,2,73,2,2,277,1,4,277,2,7,278,0,5,278,1,2,283,0,5,283,1,7,283,2,2,
/* out0170_em-eta10-phi8*/	6,50,0,3,61,1,1,61,2,9,269,1,8,277,2,7,278,0,1,
/* out0171_em-eta11-phi8*/	9,49,1,3,50,0,8,135,1,6,139,0,3,139,1,7,139,2,10,268,2,1,269,0,11,269,1,1,
/* out0172_em-eta12-phi8*/	11,38,0,2,38,1,3,49,1,1,49,2,1,50,0,1,50,2,2,134,2,1,135,0,10,135,1,3,260,1,9,269,0,2,
/* out0173_em-eta13-phi8*/	7,38,0,5,38,1,2,127,1,8,135,0,3,260,0,4,260,1,2,260,2,4,
/* out0174_em-eta14-phi8*/	8,38,0,1,38,2,6,127,0,3,127,1,3,127,2,4,251,1,2,260,0,3,260,2,2,
/* out0175_em-eta15-phi8*/	8,26,1,4,38,2,1,119,1,1,127,0,4,127,2,2,251,1,1,251,2,5,252,0,1,
/* out0176_em-eta16-phi8*/	5,26,1,4,119,1,1,119,2,5,243,1,1,251,2,5,
/* out0177_em-eta17-phi8*/	4,26,2,4,119,2,5,243,1,5,251,2,1,
/* out0178_em-eta18-phi8*/	4,15,1,1,26,2,2,112,1,4,119,2,1,
/* out0179_em-eta19-phi8*/	1,112,1,1,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	0,
/* out0185_em-eta5-phi9*/	5,86,0,1,95,0,3,95,1,14,95,2,11,96,0,2,
/* out0186_em-eta6-phi9*/	4,85,1,14,85,2,2,86,0,9,95,2,4,
/* out0187_em-eta7-phi9*/	4,73,1,2,74,0,12,74,1,1,85,2,8,
/* out0188_em-eta8-phi9*/	9,62,0,3,62,1,3,73,1,4,73,2,3,74,0,3,74,2,3,278,1,7,283,1,1,283,2,1,
/* out0189_em-eta9-phi9*/	6,62,0,10,62,1,2,62,2,4,278,0,6,278,1,6,278,2,7,
/* out0190_em-eta10-phi9*/	9,50,0,2,50,1,7,62,0,1,62,2,4,269,1,6,269,2,3,270,0,1,278,0,4,278,2,1,
/* out0191_em-eta11-phi9*/	9,50,0,2,50,1,3,50,2,5,135,1,6,135,2,2,136,0,1,269,0,2,269,1,1,269,2,11,
/* out0192_em-eta12-phi9*/	12,38,1,3,39,0,1,50,2,6,135,0,1,135,1,1,135,2,11,260,1,1,260,2,2,261,0,3,261,1,2,269,0,1,269,2,1,
/* out0193_em-eta13-phi9*/	10,38,1,7,127,1,1,127,2,1,128,0,2,128,1,3,135,0,2,135,2,2,252,1,1,260,2,7,261,0,2,
/* out0194_em-eta14-phi9*/	7,27,0,1,38,2,6,127,2,7,128,0,3,252,0,1,252,1,6,260,2,1,
/* out0195_em-eta15-phi9*/	6,26,1,1,27,0,3,38,2,1,120,1,6,127,2,2,252,0,6,
/* out0196_em-eta16-phi9*/	8,26,1,3,27,0,2,120,0,6,120,1,1,243,1,1,243,2,2,251,2,1,252,0,2,
/* out0197_em-eta17-phi9*/	9,15,1,2,26,1,1,26,2,2,112,1,1,112,2,2,119,2,1,120,0,3,243,1,5,243,2,1,
/* out0198_em-eta18-phi9*/	4,15,1,4,112,1,5,112,2,2,243,1,1,
/* out0199_em-eta19-phi9*/	2,15,1,1,112,1,2,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	0,
/* out0205_em-eta5-phi10*/	5,86,0,1,86,1,7,87,0,1,96,0,14,96,2,14,
/* out0206_em-eta6-phi10*/	4,75,0,1,86,0,5,86,1,8,86,2,14,
/* out0207_em-eta7-phi10*/	5,74,0,1,74,1,15,74,2,3,75,0,3,86,2,1,
/* out0208_em-eta8-phi10*/	5,62,1,4,63,0,6,74,2,10,278,2,1,279,0,4,
/* out0209_em-eta9-phi10*/	8,51,0,1,62,1,7,62,2,5,63,0,2,270,1,4,278,2,7,279,0,8,279,2,4,
/* out0210_em-eta10-phi10*/	5,50,1,2,51,0,9,62,2,3,270,0,7,270,1,9,
/* out0211_em-eta11-phi10*/	10,39,0,1,39,1,1,50,1,4,50,2,2,51,0,3,51,2,1,136,0,7,261,1,6,269,2,1,270,0,6,
/* out0212_em-eta12-phi10*/	9,39,0,8,50,2,1,128,1,4,135,2,1,136,0,5,136,2,5,261,0,3,261,1,6,261,2,2,
/* out0213_em-eta13-phi10*/	8,38,1,1,39,0,5,39,2,2,128,0,2,128,1,8,128,2,1,252,1,2,261,0,7,
/* out0214_em-eta14-phi10*/	7,27,0,3,27,1,3,38,2,1,120,1,1,128,0,8,252,1,6,252,2,2,
/* out0215_em-eta15-phi10*/	5,27,0,5,120,1,7,120,2,1,252,0,3,252,2,3,
/* out0216_em-eta16-phi10*/	7,27,0,2,27,2,2,120,0,3,120,1,1,120,2,3,243,2,3,252,0,3,
/* out0217_em-eta17-phi10*/	6,15,2,3,27,2,2,112,2,1,120,0,4,120,2,1,243,2,6,
/* out0218_em-eta18-phi10*/	4,15,1,3,15,2,2,112,2,6,243,1,2,
/* out0219_em-eta19-phi10*/	3,15,1,2,112,1,2,112,2,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	0,
/* out0225_em-eta5-phi11*/	4,87,0,11,87,1,12,87,2,3,96,2,2,
/* out0226_em-eta6-phi11*/	6,75,0,4,75,1,10,86,1,1,86,2,1,87,0,4,87,2,9,
/* out0227_em-eta7-phi11*/	4,63,1,1,75,0,8,75,1,2,75,2,12,
/* out0228_em-eta8-phi11*/	4,63,0,6,63,1,11,63,2,3,279,0,2,
/* out0229_em-eta9-phi11*/	9,51,1,5,63,0,2,63,2,9,270,1,2,270,2,1,271,0,2,271,1,4,279,0,2,279,2,12,
/* out0230_em-eta10-phi11*/	7,51,0,3,51,1,7,51,2,3,262,1,1,270,1,1,270,2,12,271,0,2,
/* out0231_em-eta11-phi11*/	10,39,1,3,51,2,8,136,0,3,136,2,2,261,1,2,261,2,1,262,0,2,262,1,3,270,0,2,270,2,3,
/* out0232_em-eta12-phi11*/	10,39,0,1,39,1,8,39,2,1,128,1,1,128,2,1,129,0,2,129,1,4,136,2,9,261,2,9,262,0,2,
/* out0233_em-eta13-phi11*/	8,39,2,8,128,2,9,129,0,2,252,1,1,253,0,1,253,1,4,261,0,1,261,2,4,
/* out0234_em-eta14-phi11*/	7,27,1,5,39,2,1,121,1,4,128,0,1,128,2,5,252,2,5,253,0,3,
/* out0235_em-eta15-phi11*/	6,27,1,4,27,2,2,120,2,4,121,0,4,244,1,1,252,2,5,
/* out0236_em-eta16-phi11*/	6,27,2,5,113,1,1,120,2,5,244,0,1,244,1,3,252,2,1,
/* out0237_em-eta17-phi11*/	7,15,2,3,27,2,2,113,0,1,113,1,3,120,2,2,243,2,3,244,0,3,
/* out0238_em-eta18-phi11*/	5,15,2,4,112,2,2,113,0,3,243,1,1,243,2,1,
/* out0239_em-eta19-phi11*/	3,15,1,2,112,1,1,112,2,2,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	0,
/* out0245_em-eta5-phi12*/	6,76,0,1,76,1,4,87,1,4,87,2,2,88,0,15,88,2,8,
/* out0246_em-eta6-phi12*/	5,75,1,2,76,0,15,76,1,4,76,2,5,87,2,2,
/* out0247_em-eta7-phi12*/	5,64,0,9,64,1,6,75,1,2,75,2,4,76,2,2,
/* out0248_em-eta8-phi12*/	7,52,0,1,52,1,2,63,1,4,63,2,2,64,0,7,64,2,4,271,1,2,
/* out0249_em-eta9-phi12*/	7,51,1,1,52,0,12,52,1,1,63,2,2,271,0,3,271,1,10,271,2,6,
/* out0250_em-eta10-phi12*/	9,40,0,1,40,1,2,51,1,3,51,2,2,52,0,3,52,2,2,262,1,6,271,0,9,271,2,1,
/* out0251_em-eta11-phi12*/	6,40,0,9,51,2,2,129,1,4,262,0,4,262,1,6,262,2,3,
/* out0252_em-eta12-phi12*/	10,28,1,1,39,1,4,39,2,1,40,0,4,40,2,1,129,0,2,129,1,8,129,2,3,253,1,3,262,0,7,
/* out0253_em-eta13-phi12*/	7,28,0,5,39,2,3,121,1,2,129,0,9,253,0,1,253,1,8,253,2,1,
/* out0254_em-eta14-phi12*/	5,27,1,1,28,0,5,121,1,9,121,2,1,253,0,8,
/* out0255_em-eta15-phi12*/	7,27,1,3,27,2,1,28,0,1,121,0,7,121,2,1,244,1,5,253,0,1,
/* out0256_em-eta16-phi12*/	6,16,0,2,27,2,2,113,1,4,121,0,3,244,0,1,244,1,4,
/* out0257_em-eta17-phi12*/	4,16,0,3,113,0,1,113,1,5,244,0,5,
/* out0258_em-eta18-phi12*/	4,15,2,3,16,0,1,113,0,5,244,0,2,
/* out0259_em-eta19-phi12*/	3,15,1,1,15,2,1,113,0,2,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	0,
/* out0265_em-eta5-phi13*/	6,76,1,2,77,0,14,77,1,7,77,2,1,88,0,1,88,2,8,
/* out0266_em-eta6-phi13*/	6,65,0,6,65,1,2,76,1,6,76,2,8,77,0,2,77,2,3,
/* out0267_em-eta7-phi13*/	5,64,1,10,64,2,3,65,0,8,65,2,1,76,2,1,
/* out0268_em-eta8-phi13*/	4,52,1,4,53,0,7,64,2,9,272,0,5,
/* out0269_em-eta9-phi13*/	6,52,1,9,52,2,7,263,1,4,271,2,7,272,0,8,272,2,4,
/* out0270_em-eta10-phi13*/	7,40,1,6,41,0,1,52,2,6,262,2,1,263,0,5,263,1,7,271,2,2,
/* out0271_em-eta11-phi13*/	8,40,0,2,40,1,6,40,2,3,129,2,1,130,0,6,254,1,2,262,2,9,263,0,3,
/* out0272_em-eta12-phi13*/	12,28,1,2,40,2,7,122,1,1,129,2,8,130,0,5,130,2,1,253,1,1,253,2,1,254,0,2,254,1,4,262,0,1,262,2,3,
/* out0273_em-eta13-phi13*/	9,28,0,2,28,1,6,121,1,1,122,0,2,122,1,4,129,0,1,129,2,4,253,2,8,254,0,1,
/* out0274_em-eta14-phi13*/	7,28,0,3,28,2,3,121,2,8,122,0,1,245,1,1,253,0,2,253,2,5,
/* out0275_em-eta15-phi13*/	8,16,1,2,28,2,3,114,1,1,121,0,1,121,2,6,244,1,3,244,2,3,245,0,1,
/* out0276_em-eta16-phi13*/	7,16,0,3,16,1,2,113,1,2,113,2,2,114,0,1,121,0,1,244,2,5,
/* out0277_em-eta17-phi13*/	5,16,0,4,113,1,1,113,2,5,244,0,2,244,2,2,
/* out0278_em-eta18-phi13*/	5,16,0,2,16,2,1,113,0,2,113,2,3,244,0,2,
/* out0279_em-eta19-phi13*/	3,16,0,1,16,2,1,113,0,2,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	0,
/* out0285_em-eta5-phi14*/	7,66,0,5,66,1,2,77,1,9,77,2,8,78,0,14,78,1,13,78,2,12,
/* out0286_em-eta6-phi14*/	5,65,0,1,65,1,14,65,2,2,66,0,8,77,2,4,
/* out0287_em-eta7-phi14*/	4,53,1,7,54,0,2,65,0,1,65,2,13,
/* out0288_em-eta8-phi14*/	6,53,0,7,53,1,7,53,2,6,264,0,4,272,0,3,272,2,4,
/* out0289_em-eta9-phi14*/	10,41,0,3,41,1,6,52,2,1,53,0,2,53,2,4,263,1,3,263,2,3,264,0,9,264,2,3,272,2,8,
/* out0290_em-eta10-phi14*/	6,41,0,11,41,1,1,41,2,2,263,0,4,263,1,2,263,2,10,
/* out0291_em-eta11-phi14*/	12,29,0,2,29,1,1,40,1,2,40,2,3,41,0,1,41,2,1,130,0,5,130,2,5,254,1,7,254,2,2,263,0,4,263,2,1,
/* out0292_em-eta12-phi14*/	9,28,1,1,29,0,7,40,2,2,122,1,6,122,2,1,130,2,8,254,0,5,254,1,3,254,2,2,
/* out0293_em-eta13-phi14*/	9,28,1,6,28,2,1,29,0,1,122,0,4,122,1,5,122,2,3,245,1,3,253,2,1,254,0,6,
/* out0294_em-eta14-phi14*/	4,28,2,6,114,1,2,122,0,7,245,1,7,
/* out0295_em-eta15-phi14*/	6,16,1,3,17,0,1,28,2,2,114,1,8,244,2,1,245,0,6,
/* out0296_em-eta16-phi14*/	6,16,1,5,114,0,6,114,1,1,237,1,1,244,2,3,245,0,1,
/* out0297_em-eta17-phi14*/	7,16,1,1,16,2,3,107,1,1,113,2,4,114,0,1,237,1,2,244,2,2,
/* out0298_em-eta18-phi14*/	4,16,2,3,107,1,2,113,2,2,237,1,1,
/* out0299_em-eta19-phi14*/	2,16,2,1,107,1,2,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	0,
/* out0305_em-eta5-phi15*/	8,66,1,14,66,2,2,67,0,16,67,1,10,67,2,1,78,0,2,78,1,3,78,2,4,
/* out0306_em-eta6-phi15*/	5,54,0,1,54,1,8,55,0,2,66,0,3,66,2,14,
/* out0307_em-eta7-phi15*/	3,54,0,12,54,1,5,54,2,6,
/* out0308_em-eta8-phi15*/	7,42,0,6,42,1,4,53,1,2,53,2,5,54,0,1,54,2,2,264,1,4,
/* out0309_em-eta9-phi15*/	6,41,1,8,42,0,7,53,2,1,264,0,3,264,1,7,264,2,11,
/* out0310_em-eta10-phi15*/	6,30,0,1,41,1,1,41,2,11,255,1,13,263,2,2,264,2,2,
/* out0311_em-eta11-phi15*/	8,29,1,9,41,2,2,123,0,9,123,1,4,130,2,2,254,2,3,255,0,9,255,1,1,
/* out0312_em-eta12-phi15*/	8,29,0,4,29,1,2,29,2,4,122,2,2,123,0,7,123,2,9,246,1,3,254,2,8,
/* out0313_em-eta13-phi15*/	12,17,1,2,29,0,2,29,2,3,115,1,2,122,2,8,123,2,1,245,1,3,245,2,2,246,0,1,246,1,1,254,0,2,254,2,1,
/* out0314_em-eta14-phi15*/	11,17,0,5,17,1,1,28,2,1,114,1,2,114,2,2,115,0,1,115,1,2,122,0,2,122,2,2,245,1,2,245,2,5,
/* out0315_em-eta15-phi15*/	5,17,0,5,114,1,2,114,2,5,245,0,6,245,2,1,
/* out0316_em-eta16-phi15*/	7,16,1,3,17,0,1,114,0,5,114,2,2,237,1,1,237,2,4,245,0,1,
/* out0317_em-eta17-phi15*/	4,16,2,4,107,2,4,114,0,2,237,1,4,
/* out0318_em-eta18-phi15*/	4,16,2,3,107,1,3,107,2,1,237,1,2,
/* out0319_em-eta19-phi15*/	1,107,1,3,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	0,
/* out0325_em-eta5-phi16*/	6,55,0,1,55,1,10,56,0,5,56,1,6,67,1,6,67,2,15,
/* out0326_em-eta6-phi16*/	5,43,1,1,54,1,1,55,0,13,55,1,4,55,2,10,
/* out0327_em-eta7-phi16*/	4,43,0,10,43,1,3,54,1,2,54,2,8,
/* out0328_em-eta8-phi16*/	5,42,0,1,42,1,12,42,2,4,43,0,2,264,1,1,
/* out0329_em-eta9-phi16*/	7,30,1,4,42,0,2,42,2,10,256,0,16,256,1,3,256,2,4,264,1,4,
/* out0330_em-eta10-phi16*/	5,30,0,9,30,1,4,255,1,2,255,2,12,256,2,3,
/* out0331_em-eta11-phi16*/	7,29,1,4,30,0,6,30,2,1,123,1,6,246,1,2,255,0,7,255,2,4,
/* out0332_em-eta12-phi16*/	8,18,0,2,29,2,7,115,1,1,123,1,6,123,2,6,246,0,1,246,1,9,246,2,1,
/* out0333_em-eta13-phi16*/	8,17,1,5,18,0,1,29,2,2,115,1,10,115,2,1,245,2,1,246,0,8,246,1,1,
/* out0334_em-eta14-phi16*/	8,17,0,1,17,1,4,17,2,1,115,0,8,115,1,1,238,1,2,245,2,5,246,0,1,
/* out0335_em-eta15-phi16*/	9,17,0,2,17,2,3,108,1,2,114,2,4,115,0,2,238,0,1,238,1,2,245,0,1,245,2,2,
/* out0336_em-eta16-phi16*/	7,7,2,1,17,0,1,17,2,2,108,1,3,114,0,1,114,2,3,237,2,6,
/* out0337_em-eta17-phi16*/	6,7,1,3,107,2,5,108,0,1,237,0,2,237,1,1,237,2,2,
/* out0338_em-eta18-phi16*/	5,7,1,3,107,0,2,107,1,1,107,2,3,237,1,3,
/* out0339_em-eta19-phi16*/	1,107,1,3,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	0,
/* out0345_em-eta5-phi17*/	5,44,1,5,55,1,1,56,0,11,56,1,10,56,2,16,
/* out0346_em-eta6-phi17*/	5,43,1,3,44,0,15,44,1,3,55,1,1,55,2,6,
/* out0347_em-eta7-phi17*/	4,43,0,2,43,1,9,43,2,11,44,0,1,
/* out0348_em-eta8-phi17*/	5,31,0,4,31,1,8,42,2,1,43,0,2,43,2,5,
/* out0349_em-eta9-phi17*/	5,30,1,3,31,0,12,42,2,1,256,1,13,256,2,4,
/* out0350_em-eta10-phi17*/	4,30,1,5,30,2,9,247,1,11,256,2,5,
/* out0351_em-eta11-phi17*/	7,18,1,5,30,2,6,116,0,3,116,1,3,246,2,1,247,0,7,247,1,5,
/* out0352_em-eta12-phi17*/	8,18,0,7,18,1,3,115,2,1,116,0,13,116,1,1,116,2,7,246,2,11,247,0,1,
/* out0353_em-eta13-phi17*/	7,17,1,2,18,0,6,115,2,10,116,2,1,238,1,1,246,0,5,246,2,3,
/* out0354_em-eta14-phi17*/	6,17,1,2,17,2,4,108,1,1,115,0,5,115,2,4,238,1,8,
/* out0355_em-eta15-phi17*/	4,17,2,5,108,1,7,238,0,4,238,1,3,
/* out0356_em-eta16-phi17*/	6,7,2,4,17,2,1,108,0,3,108,1,3,237,2,3,238,0,3,
/* out0357_em-eta17-phi17*/	6,7,1,2,7,2,2,107,2,2,108,0,4,237,0,9,237,2,1,
/* out0358_em-eta18-phi17*/	5,7,1,3,107,0,8,107,2,1,237,0,5,237,1,1,
/* out0359_em-eta19-phi17*/	2,107,0,6,107,1,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	0,
/* out0365_em-eta5-phi18*/	5,33,1,1,44,1,5,45,0,16,45,1,15,45,2,9,
/* out0366_em-eta6-phi18*/	5,32,1,3,33,0,6,33,1,1,44,1,3,44,2,15,
/* out0367_em-eta7-phi18*/	4,32,0,11,32,1,9,32,2,2,44,2,1,
/* out0368_em-eta8-phi18*/	5,20,0,1,31,1,8,31,2,4,32,0,5,32,2,2,
/* out0369_em-eta9-phi18*/	6,19,1,3,20,0,1,31,2,12,248,0,16,248,1,6,248,2,5,
/* out0370_em-eta10-phi18*/	4,19,0,9,19,1,5,247,2,11,248,2,5,
/* out0371_em-eta11-phi18*/	7,18,1,5,19,0,6,110,0,1,116,1,5,239,1,1,247,0,7,247,2,5,
/* out0372_em-eta12-phi18*/	7,18,1,3,18,2,7,109,1,1,116,1,7,116,2,6,239,1,11,247,0,1,
/* out0373_em-eta13-phi18*/	7,8,1,2,18,2,6,109,1,10,116,2,2,238,2,1,239,0,5,239,1,3,
/* out0374_em-eta14-phi18*/	6,8,0,4,8,1,2,108,2,1,109,0,5,109,1,4,238,2,8,
/* out0375_em-eta15-phi18*/	4,8,0,5,108,2,7,238,0,4,238,2,3,
/* out0376_em-eta16-phi18*/	6,7,2,4,8,0,1,108,0,3,108,2,3,232,2,3,238,0,3,
/* out0377_em-eta17-phi18*/	6,7,0,2,7,1,1,7,2,3,103,2,2,108,0,4,232,1,4,
/* out0378_em-eta18-phi18*/	4,7,1,3,103,1,3,103,2,1,232,1,3,
/* out0379_em-eta19-phi18*/	1,103,1,3,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	0,
/* out0385_em-eta5-phi19*/	7,33,1,10,33,2,1,34,0,16,34,1,12,34,2,2,45,1,1,45,2,7,
/* out0386_em-eta6-phi19*/	5,21,1,1,32,1,1,33,0,10,33,1,4,33,2,13,
/* out0387_em-eta7-phi19*/	4,21,0,8,21,1,2,32,1,3,32,2,10,
/* out0388_em-eta8-phi19*/	6,20,0,4,20,1,12,20,2,1,32,2,2,241,1,1,248,1,1,
/* out0389_em-eta9-phi19*/	7,19,1,4,20,0,10,20,2,2,241,0,10,241,2,1,248,1,9,248,2,3,
/* out0390_em-eta10-phi19*/	5,19,1,4,19,2,9,240,1,12,240,2,2,248,2,3,
/* out0391_em-eta11-phi19*/	8,9,1,4,19,0,1,19,2,6,110,0,3,110,1,5,239,2,2,240,0,7,240,1,4,
/* out0392_em-eta12-phi19*/	9,9,0,7,18,2,2,109,2,1,110,0,12,110,1,1,110,2,7,239,0,1,239,1,1,239,2,9,
/* out0393_em-eta13-phi19*/	8,8,1,5,9,0,2,18,2,1,109,1,1,109,2,10,233,1,1,239,0,8,239,2,1,
/* out0394_em-eta14-phi19*/	8,8,0,1,8,1,4,8,2,1,109,0,8,109,2,1,233,1,5,238,2,2,239,0,1,
/* out0395_em-eta15-phi19*/	9,8,0,3,8,2,2,104,1,4,108,2,2,109,0,2,233,0,1,233,1,2,238,0,1,238,2,2,
/* out0396_em-eta16-phi19*/	8,7,0,1,7,2,2,8,0,2,8,2,1,104,0,1,104,1,3,108,2,3,232,2,6,
/* out0397_em-eta17-phi19*/	5,7,0,8,103,2,5,108,0,1,232,1,2,232,2,2,
/* out0398_em-eta18-phi19*/	5,7,0,4,7,1,1,103,1,2,103,2,3,232,1,3,
/* out0399_em-eta19-phi19*/	1,103,1,3,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	0,
/* out0405_em-eta5-phi20*/	7,22,0,2,22,1,14,23,0,4,23,1,3,23,2,2,34,1,4,34,2,14,
/* out0406_em-eta6-phi20*/	5,21,1,8,21,2,1,22,0,14,22,2,3,33,2,2,
/* out0407_em-eta7-phi20*/	3,21,0,6,21,1,5,21,2,12,
/* out0408_em-eta8-phi20*/	7,11,0,5,11,1,2,20,1,4,20,2,6,21,0,2,21,2,1,241,1,4,
/* out0409_em-eta9-phi20*/	6,10,1,8,11,0,1,20,2,7,241,0,6,241,1,6,241,2,11,
/* out0410_em-eta10-phi20*/	6,10,0,11,10,1,1,19,2,1,235,1,2,240,2,13,241,2,1,
/* out0411_em-eta11-phi20*/	7,9,1,9,10,0,2,106,0,2,110,1,7,234,1,3,240,0,9,240,2,1,
/* out0412_em-eta12-phi20*/	8,9,0,4,9,1,2,9,2,4,105,1,2,110,1,3,110,2,8,234,1,8,239,2,3,
/* out0413_em-eta13-phi20*/	12,8,1,2,9,0,3,9,2,2,105,1,8,109,2,2,110,2,1,233,1,2,233,2,3,234,0,2,234,1,1,239,0,1,239,2,1,
/* out0414_em-eta14-phi20*/	11,1,0,1,8,1,1,8,2,5,104,1,2,104,2,2,105,0,2,105,1,2,109,0,1,109,2,2,233,1,5,233,2,2,
/* out0415_em-eta15-phi20*/	5,8,2,5,104,1,5,104,2,2,233,0,6,233,1,1,
/* out0416_em-eta16-phi20*/	7,0,1,3,8,2,1,104,0,5,104,1,2,232,0,1,232,2,4,233,0,1,
/* out0417_em-eta17-phi20*/	6,0,0,4,103,2,4,104,0,2,232,0,6,232,1,1,232,2,1,
/* out0418_em-eta18-phi20*/	6,0,0,3,7,0,1,103,0,7,103,1,1,103,2,1,232,1,2,
/* out0419_em-eta19-phi20*/	1,103,1,3,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	0,
/* out0425_em-eta5-phi21*/	7,13,0,8,13,1,9,22,1,2,22,2,5,23,0,12,23,1,13,23,2,14,
/* out0426_em-eta6-phi21*/	5,12,0,2,12,1,14,12,2,1,13,0,4,22,2,8,
/* out0427_em-eta7-phi21*/	4,11,1,7,12,0,13,12,2,1,21,2,2,
/* out0428_em-eta8-phi21*/	5,11,0,6,11,1,7,11,2,7,236,0,7,241,1,2,
/* out0429_em-eta9-phi21*/	11,3,0,1,10,1,6,10,2,3,11,0,4,11,2,2,235,1,3,235,2,3,236,0,5,236,2,3,241,1,3,241,2,3,
/* out0430_em-eta10-phi21*/	6,10,0,2,10,1,1,10,2,11,235,0,4,235,1,10,235,2,2,
/* out0431_em-eta11-phi21*/	12,2,0,3,2,1,2,9,1,1,9,2,2,10,0,1,10,2,1,106,0,10,106,2,1,234,1,2,234,2,7,235,0,4,235,1,1,
/* out0432_em-eta12-phi21*/	10,1,1,1,2,0,2,9,2,7,105,1,1,105,2,6,106,0,2,106,2,7,234,0,5,234,1,2,234,2,3,
/* out0433_em-eta13-phi21*/	9,1,0,1,1,1,6,9,2,1,105,0,4,105,1,3,105,2,5,229,1,1,233,2,3,234,0,6,
/* out0434_em-eta14-phi21*/	4,1,0,6,104,2,2,105,0,7,233,2,7,
/* out0435_em-eta15-phi21*/	6,0,1,3,1,0,2,8,2,1,104,2,8,228,1,1,233,0,6,
/* out0436_em-eta16-phi21*/	6,0,1,5,104,0,6,104,2,1,228,1,3,232,0,2,233,0,1,
/* out0437_em-eta17-phi21*/	7,0,0,3,0,1,1,100,1,4,103,0,1,104,0,1,228,1,2,232,0,6,
/* out0438_em-eta18-phi21*/	6,0,0,3,100,1,2,103,0,6,228,0,1,232,0,1,232,1,1,
/* out0439_em-eta19-phi21*/	4,0,0,1,100,0,1,103,0,2,103,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	0,
/* out0445_em-eta5-phi22*/	6,5,1,2,6,0,8,6,2,1,13,0,1,13,1,7,13,2,14,
/* out0446_em-eta6-phi22*/	6,5,0,8,5,1,6,12,1,2,12,2,6,13,0,3,13,2,2,
/* out0447_em-eta7-phi22*/	5,4,0,3,4,1,10,5,0,1,12,0,1,12,2,8,
/* out0448_em-eta8-phi22*/	5,3,1,4,4,0,9,11,2,7,236,0,4,236,2,1,
/* out0449_em-eta9-phi22*/	5,3,0,7,3,1,9,231,1,7,235,2,4,236,2,12,
/* out0450_em-eta10-phi22*/	9,2,1,6,3,0,6,10,2,1,230,1,1,230,2,3,231,0,1,231,1,2,235,0,5,235,2,7,
/* out0451_em-eta11-phi22*/	10,2,0,3,2,1,6,2,2,2,102,1,1,102,2,3,106,0,2,106,2,3,230,1,9,234,2,2,235,0,3,
/* out0452_em-eta12-phi22*/	11,1,1,2,2,0,7,102,1,8,105,2,1,106,2,5,229,1,1,229,2,1,230,0,1,230,1,3,234,0,2,234,2,4,
/* out0453_em-eta13-phi22*/	10,1,1,6,1,2,2,101,2,1,102,0,1,102,1,4,105,0,2,105,2,4,229,1,8,229,2,3,234,0,1,
/* out0454_em-eta14-phi22*/	8,1,0,3,1,2,3,101,1,8,101,2,1,105,0,1,229,0,2,229,1,5,233,2,1,
/* out0455_em-eta15-phi22*/	9,0,1,2,1,0,3,101,0,2,101,1,6,104,2,1,228,1,3,228,2,3,229,0,1,233,0,1,
/* out0456_em-eta16-phi22*/	9,0,1,2,0,2,3,100,1,2,100,2,3,101,0,2,104,0,1,228,0,1,228,1,5,228,2,1,
/* out0457_em-eta17-phi22*/	6,0,2,4,100,0,1,100,1,5,100,2,1,228,0,3,228,1,2,
/* out0458_em-eta18-phi22*/	5,0,0,1,0,2,2,100,0,2,100,1,3,228,0,2,
/* out0459_em-eta19-phi22*/	3,0,0,1,0,2,1,100,0,3,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	0,
/* out0465_em-eta5-phi23*/	4,5,1,4,5,2,1,6,0,8,6,2,15,
/* out0466_em-eta6-phi23*/	3,5,0,5,5,1,4,5,2,15,
/* out0467_em-eta7-phi23*/	3,4,1,6,4,2,9,5,0,2,
/* out0468_em-eta8-phi23*/	5,3,1,2,3,2,1,4,0,4,4,2,7,231,2,2,
/* out0469_em-eta9-phi23*/	5,3,1,1,3,2,12,231,0,3,231,1,6,231,2,14,
/* out0470_em-eta10-phi23*/	7,2,1,2,2,2,1,3,0,2,3,2,3,230,2,6,231,0,12,231,1,1,
/* out0471_em-eta11-phi23*/	5,2,2,9,102,2,4,230,0,4,230,1,3,230,2,7,
/* out0472_em-eta12-phi23*/	8,1,1,1,2,0,1,2,2,4,102,0,6,102,1,3,102,2,9,229,2,4,230,0,11,
/* out0473_em-eta13-phi23*/	6,1,2,5,101,2,2,102,0,9,229,0,1,229,1,1,229,2,8,
/* out0474_em-eta14-phi23*/	5,1,2,5,101,0,1,101,1,1,101,2,9,229,0,8,
/* out0475_em-eta15-phi23*/	6,1,2,1,101,0,8,101,1,1,101,2,3,228,2,8,229,0,4,
/* out0476_em-eta16-phi23*/	5,0,2,2,100,2,7,101,0,3,228,0,2,228,2,4,
/* out0477_em-eta17-phi23*/	4,0,2,3,100,0,1,100,2,5,228,0,5,
/* out0478_em-eta18-phi23*/	3,0,2,1,100,0,5,228,0,2,
/* out0479_em-eta19-phi23*/	1,100,0,3
};