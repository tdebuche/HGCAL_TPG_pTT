parameter integer matrixH [0:6353] = {
/* num inputs = 251(in0-in250) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 10 */
//* total number of input in adders 1957 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	1,99,0,13,
/* out0002_em-eta2-phi0*/	2,99,0,3,99,1,14,
/* out0003_em-eta3-phi0*/	2,98,0,16,99,1,2,
/* out0004_em-eta4-phi0*/	2,87,2,2,98,1,16,
/* out0005_em-eta5-phi0*/	6,86,0,3,86,1,6,87,1,8,87,2,13,97,0,16,97,1,2,
/* out0006_em-eta6-phi0*/	6,85,1,1,86,0,13,86,1,2,86,2,7,96,0,2,97,1,14,
/* out0007_em-eta7-phi0*/	5,85,0,13,85,1,4,85,2,1,96,0,14,96,1,4,
/* out0008_em-eta8-phi0*/	6,84,0,3,84,1,3,85,0,3,85,2,3,96,1,12,96,2,4,
/* out0009_em-eta9-phi0*/	4,84,0,12,84,2,1,95,0,3,96,2,12,
/* out0010_em-eta10-phi0*/	6,83,0,3,83,1,1,84,0,1,84,2,1,95,0,13,95,1,3,
/* out0011_em-eta11-phi0*/	4,83,0,9,104,0,2,104,1,6,95,1,13,
/* out0012_em-eta12-phi0*/	6,82,0,1,82,1,1,83,0,2,104,0,7,104,1,3,104,2,4,
/* out0013_em-eta13-phi0*/	5,82,0,6,103,0,1,103,1,4,104,0,7,104,2,5,
/* out0014_em-eta14-phi0*/	4,82,0,4,103,0,6,103,1,3,103,2,1,
/* out0015_em-eta15-phi0*/	3,81,0,1,103,0,3,103,2,5,
/* out0016_em-eta16-phi0*/	4,81,0,3,102,0,2,102,1,4,103,0,6,
/* out0017_em-eta17-phi0*/	3,81,0,3,102,0,5,102,1,1,
/* out0018_em-eta18-phi0*/	2,102,0,8,102,2,2,
/* out0019_em-eta19-phi0*/	2,102,0,1,102,2,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	1,99,3,13,
/* out0022_em-eta2-phi1*/	2,99,2,14,99,3,3,
/* out0023_em-eta3-phi1*/	2,98,3,16,99,2,2,
/* out0024_em-eta4-phi1*/	4,80,1,3,87,1,1,87,2,1,98,2,16,
/* out0025_em-eta5-phi1*/	7,80,0,16,80,1,4,80,2,3,86,1,5,87,1,7,97,2,2,97,3,16,
/* out0026_em-eta6-phi1*/	8,79,0,10,79,1,2,80,2,1,85,1,1,86,1,3,86,2,9,96,5,2,97,2,14,
/* out0027_em-eta7-phi1*/	6,78,0,2,79,0,4,85,1,10,85,2,7,96,4,4,96,5,14,
/* out0028_em-eta8-phi1*/	5,78,0,6,84,1,8,85,2,5,96,3,4,96,4,12,
/* out0029_em-eta9-phi1*/	4,84,1,5,84,2,10,95,3,3,96,3,12,
/* out0030_em-eta10-phi1*/	5,77,0,1,83,1,9,84,2,3,95,2,3,95,3,13,
/* out0031_em-eta11-phi1*/	6,83,0,2,83,1,3,83,2,6,100,2,9,104,1,3,95,2,13,
/* out0032_em-eta12-phi1*/	6,82,1,4,83,2,5,98,0,3,100,2,1,104,1,4,104,2,5,
/* out0033_em-eta13-phi1*/	6,82,0,3,82,1,4,82,2,1,98,0,6,103,1,3,104,2,2,
/* out0034_em-eta14-phi1*/	4,82,0,2,82,2,4,103,1,6,103,2,3,
/* out0035_em-eta15-phi1*/	5,81,0,1,81,1,3,82,2,2,97,0,1,103,2,6,
/* out0036_em-eta16-phi1*/	4,81,0,3,81,1,1,97,0,1,102,1,6,
/* out0037_em-eta17-phi1*/	3,81,0,3,102,1,3,102,2,3,
/* out0038_em-eta18-phi1*/	3,81,0,2,81,2,1,102,2,5,
/* out0039_em-eta19-phi1*/	1,102,2,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	1,104,0,13,
/* out0042_em-eta2-phi2*/	2,104,0,3,104,1,14,
/* out0043_em-eta3-phi2*/	2,103,0,16,104,1,2,
/* out0044_em-eta4-phi2*/	2,80,1,2,103,1,16,
/* out0045_em-eta5-phi2*/	6,74,0,8,74,1,2,80,1,7,80,2,11,102,0,16,102,1,2,
/* out0046_em-eta6-phi2*/	7,74,0,4,79,0,2,79,1,14,79,2,7,80,2,1,101,0,2,102,1,14,
/* out0047_em-eta7-phi2*/	6,73,0,2,78,0,1,78,1,11,79,2,9,101,0,14,101,1,4,
/* out0048_em-eta8-phi2*/	5,78,0,7,78,1,2,78,2,9,101,1,12,101,2,4,
/* out0049_em-eta9-phi2*/	6,77,0,6,77,1,7,78,2,1,84,2,1,100,0,3,101,2,12,
/* out0050_em-eta10-phi2*/	5,77,0,9,77,2,3,83,1,2,100,0,13,100,1,3,
/* out0051_em-eta11-phi2*/	7,76,0,4,76,1,1,83,1,1,83,2,4,100,1,10,100,2,6,100,1,13,
/* out0052_em-eta12-phi2*/	6,76,0,6,82,1,2,83,2,1,98,0,1,98,1,9,100,1,4,
/* out0053_em-eta13-phi2*/	5,82,1,5,82,2,2,98,0,5,98,1,1,98,2,5,
/* out0054_em-eta14-phi2*/	7,75,0,1,82,2,6,97,0,1,97,1,3,98,0,1,98,2,3,103,2,1,
/* out0055_em-eta15-phi2*/	4,81,1,4,82,2,1,97,0,7,97,1,1,
/* out0056_em-eta16-phi2*/	3,81,1,4,97,0,5,102,1,1,
/* out0057_em-eta17-phi2*/	4,81,2,4,96,1,1,102,1,1,102,2,2,
/* out0058_em-eta18-phi2*/	3,81,2,3,96,1,3,102,2,2,
/* out0059_em-eta19-phi2*/	1,96,0,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	1,104,3,13,
/* out0062_em-eta2-phi3*/	2,104,2,14,104,3,3,
/* out0063_em-eta3-phi3*/	2,103,3,16,104,2,2,
/* out0064_em-eta4-phi3*/	3,69,0,3,69,2,7,103,2,16,
/* out0065_em-eta5-phi3*/	9,68,0,1,69,0,1,69,1,8,69,2,9,74,0,2,74,1,14,74,2,7,102,2,2,102,3,16,
/* out0066_em-eta6-phi3*/	7,68,0,2,73,0,3,73,1,12,74,0,2,74,2,9,101,5,2,102,2,14,
/* out0067_em-eta7-phi3*/	7,72,1,1,73,0,11,73,1,1,73,2,8,78,1,2,101,4,4,101,5,14,
/* out0068_em-eta8-phi3*/	6,72,0,10,72,1,3,78,1,1,78,2,6,101,3,4,101,4,12,
/* out0069_em-eta9-phi3*/	5,72,0,4,77,1,9,77,2,3,100,3,3,101,3,12,
/* out0070_em-eta10-phi3*/	5,71,0,1,76,1,1,77,2,10,100,2,3,100,3,13,
/* out0071_em-eta11-phi3*/	6,76,0,1,76,1,10,100,1,2,101,0,8,101,2,9,100,2,13,
/* out0072_em-eta12-phi3*/	5,76,0,4,76,2,5,98,1,5,101,1,2,101,2,7,
/* out0073_em-eta13-phi3*/	7,75,0,1,75,1,3,76,0,1,76,2,2,98,1,1,98,2,7,99,1,3,
/* out0074_em-eta14-phi3*/	4,75,0,6,97,1,6,98,2,1,99,1,2,
/* out0075_em-eta15-phi3*/	5,75,0,4,81,1,1,97,0,1,97,1,4,97,2,3,
/* out0076_em-eta16-phi3*/	3,81,1,3,81,2,2,97,2,6,
/* out0077_em-eta17-phi3*/	2,81,2,4,96,1,5,
/* out0078_em-eta18-phi3*/	3,81,2,2,96,0,2,96,1,3,
/* out0079_em-eta19-phi3*/	1,96,0,3,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	1,109,0,13,
/* out0082_em-eta2-phi4*/	2,109,0,3,109,1,14,
/* out0083_em-eta3-phi4*/	2,108,0,16,109,1,2,
/* out0084_em-eta4-phi4*/	2,69,0,3,108,1,16,
/* out0085_em-eta5-phi4*/	9,68,0,3,68,1,14,68,2,1,69,0,9,69,1,8,70,0,5,70,1,6,107,0,16,107,1,2,
/* out0086_em-eta6-phi4*/	7,67,1,3,68,0,10,68,2,9,73,1,3,73,2,1,106,0,2,107,1,14,
/* out0087_em-eta7-phi4*/	6,67,0,12,67,1,1,72,1,3,73,2,7,106,0,14,106,1,4,
/* out0088_em-eta8-phi4*/	5,72,0,1,72,1,9,72,2,8,106,1,12,106,2,4,
/* out0089_em-eta9-phi4*/	6,71,0,1,71,1,7,72,0,1,72,2,7,105,0,3,106,2,12,
/* out0090_em-eta10-phi4*/	5,71,0,11,71,1,1,71,2,1,105,0,13,105,1,3,
/* out0091_em-eta11-phi4*/	8,56,1,1,71,0,3,71,2,1,76,1,4,76,2,2,101,0,8,101,1,6,105,1,13,
/* out0092_em-eta12-phi4*/	4,56,1,2,76,2,6,99,2,5,101,1,8,
/* out0093_em-eta13-phi4*/	5,75,1,7,76,2,1,99,0,1,99,1,5,99,2,5,
/* out0094_em-eta14-phi4*/	6,75,0,2,75,1,2,75,2,2,97,1,1,99,0,2,99,1,6,
/* out0095_em-eta15-phi4*/	5,75,0,2,75,2,4,92,1,2,97,1,1,97,2,4,
/* out0096_em-eta16-phi4*/	6,75,2,1,88,1,2,92,1,2,96,1,1,96,2,1,97,2,3,
/* out0097_em-eta17-phi4*/	3,88,1,3,96,1,2,96,2,3,
/* out0098_em-eta18-phi4*/	5,88,0,2,88,1,1,96,0,3,96,1,1,96,2,2,
/* out0099_em-eta19-phi4*/	1,96,0,4,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	1,109,3,13,
/* out0102_em-eta2-phi5*/	2,109,2,14,109,3,3,
/* out0103_em-eta3-phi5*/	2,108,3,16,109,2,2,
/* out0104_em-eta4-phi5*/	1,108,2,16,
/* out0105_em-eta5-phi5*/	9,63,0,2,63,1,7,68,1,2,68,2,2,70,0,11,70,1,10,70,2,16,107,2,2,107,3,16,
/* out0106_em-eta6-phi5*/	5,63,0,14,67,1,8,68,2,4,106,5,2,107,2,14,
/* out0107_em-eta7-phi5*/	5,67,0,3,67,1,4,67,2,15,106,4,4,106,5,14,
/* out0108_em-eta8-phi5*/	7,61,1,8,61,2,7,67,0,1,67,2,1,72,2,1,106,3,4,106,4,12,
/* out0109_em-eta9-phi5*/	4,61,1,8,71,1,6,105,3,3,106,3,12,
/* out0110_em-eta10-phi5*/	4,71,1,2,71,2,11,105,2,3,105,3,13,
/* out0111_em-eta11-phi5*/	6,56,1,1,56,2,7,71,2,3,94,0,9,94,2,5,105,2,13,
/* out0112_em-eta12-phi5*/	5,56,1,8,56,2,1,94,1,1,94,2,11,99,2,2,
/* out0113_em-eta13-phi5*/	4,56,1,4,75,1,3,99,0,7,99,2,4,
/* out0114_em-eta14-phi5*/	4,75,1,1,75,2,5,92,2,2,99,0,6,
/* out0115_em-eta15-phi5*/	4,75,2,4,88,1,1,92,1,3,92,2,5,
/* out0116_em-eta16-phi5*/	2,88,1,4,92,1,7,
/* out0117_em-eta17-phi5*/	4,88,0,1,88,1,3,92,1,2,96,2,4,
/* out0118_em-eta18-phi5*/	2,88,0,4,96,2,5,
/* out0119_em-eta19-phi5*/	2,96,0,3,96,2,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	1,114,0,13,
/* out0122_em-eta2-phi6*/	2,114,0,3,114,1,14,
/* out0123_em-eta3-phi6*/	2,113,0,16,114,1,2,
/* out0124_em-eta4-phi6*/	1,113,1,16,
/* out0125_em-eta5-phi6*/	9,63,1,8,63,2,2,64,1,2,64,2,2,65,0,11,65,1,14,65,2,16,112,0,16,112,1,2,
/* out0126_em-eta6-phi6*/	6,62,2,8,63,1,1,63,2,14,64,1,4,111,0,2,112,1,14,
/* out0127_em-eta7-phi6*/	6,61,2,1,62,0,3,62,1,15,62,2,4,111,0,14,111,1,4,
/* out0128_em-eta8-phi6*/	7,58,1,1,61,0,8,61,2,8,62,0,1,62,1,1,111,1,12,111,2,4,
/* out0129_em-eta9-phi6*/	4,57,2,6,61,0,8,110,0,3,111,2,12,
/* out0130_em-eta10-phi6*/	4,57,1,11,57,2,2,110,0,13,110,1,3,
/* out0131_em-eta11-phi6*/	6,56,0,1,56,2,7,57,1,3,94,0,7,94,1,5,110,1,13,
/* out0132_em-eta12-phi6*/	4,56,0,8,56,2,1,93,2,2,94,1,10,
/* out0133_em-eta13-phi6*/	4,56,0,4,89,2,3,93,1,7,93,2,4,
/* out0134_em-eta14-phi6*/	4,89,1,5,89,2,1,92,2,3,93,1,6,
/* out0135_em-eta15-phi6*/	4,88,2,1,89,1,4,92,0,3,92,2,5,
/* out0136_em-eta16-phi6*/	3,88,1,1,88,2,4,92,0,6,
/* out0137_em-eta17-phi6*/	5,88,0,2,88,1,1,88,2,2,92,0,2,105,1,3,
/* out0138_em-eta18-phi6*/	2,88,0,4,105,1,4,
/* out0139_em-eta19-phi6*/	2,105,0,2,105,1,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	1,114,3,13,
/* out0142_em-eta2-phi7*/	2,114,2,14,114,3,3,
/* out0143_em-eta3-phi7*/	2,113,3,16,114,2,2,
/* out0144_em-eta4-phi7*/	2,66,1,3,113,2,16,
/* out0145_em-eta5-phi7*/	10,64,0,3,64,1,1,64,2,14,65,0,5,65,1,2,66,0,16,66,1,9,66,2,2,112,2,2,112,3,16,
/* out0146_em-eta6-phi7*/	7,59,1,1,59,2,3,62,2,3,64,0,10,64,1,9,111,5,2,112,2,14,
/* out0147_em-eta7-phi7*/	6,58,2,3,59,1,7,62,0,12,62,2,1,111,4,4,111,5,14,
/* out0148_em-eta8-phi7*/	5,58,0,1,58,1,8,58,2,9,111,3,4,111,4,12,
/* out0149_em-eta9-phi7*/	6,57,0,1,57,2,7,58,0,1,58,1,7,110,3,3,111,3,12,
/* out0150_em-eta10-phi7*/	5,57,0,11,57,1,1,57,2,1,110,2,3,110,3,13,
/* out0151_em-eta11-phi7*/	9,56,0,1,57,0,3,57,1,1,90,1,2,90,2,4,95,0,10,95,1,1,95,2,5,110,2,13,
/* out0152_em-eta12-phi7*/	4,56,0,2,90,1,6,93,2,5,95,2,10,
/* out0153_em-eta13-phi7*/	5,89,2,7,90,1,1,93,0,5,93,1,1,93,2,5,
/* out0154_em-eta14-phi7*/	6,89,0,2,89,1,2,89,2,2,93,0,6,93,1,2,106,2,1,
/* out0155_em-eta15-phi7*/	6,89,0,2,89,1,4,92,0,2,92,2,1,106,1,4,106,2,1,
/* out0156_em-eta16-phi7*/	6,88,2,4,89,1,1,92,0,3,105,1,1,105,2,1,106,1,3,
/* out0157_em-eta17-phi7*/	3,88,2,4,105,1,4,105,2,1,
/* out0158_em-eta18-phi7*/	4,88,0,3,88,2,1,105,0,2,105,1,3,
/* out0159_em-eta19-phi7*/	1,105,0,4,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	1,119,0,13,
/* out0162_em-eta2-phi8*/	2,119,0,3,119,1,14,
/* out0163_em-eta3-phi8*/	2,118,0,16,119,1,2,
/* out0164_em-eta4-phi8*/	3,66,1,3,66,2,3,118,1,16,
/* out0165_em-eta5-phi8*/	8,60,0,2,60,1,7,60,2,14,64,0,1,66,1,1,66,2,11,117,0,16,117,1,2,
/* out0166_em-eta6-phi8*/	7,59,0,3,59,2,12,60,0,2,60,1,9,64,0,2,116,0,2,117,1,14,
/* out0167_em-eta7-phi8*/	7,58,2,1,59,0,11,59,1,8,59,2,1,92,2,2,116,0,14,116,1,4,
/* out0168_em-eta8-phi8*/	6,58,0,10,58,2,3,92,1,6,92,2,1,116,1,12,116,2,4,
/* out0169_em-eta9-phi8*/	5,58,0,4,91,1,3,91,2,9,115,0,3,116,2,12,
/* out0170_em-eta10-phi8*/	5,57,0,1,90,2,1,91,1,10,115,0,13,115,1,3,
/* out0171_em-eta11-phi8*/	6,90,0,1,90,2,10,95,0,6,95,1,8,108,1,2,115,1,13,
/* out0172_em-eta12-phi8*/	5,90,0,4,90,1,5,95,1,7,95,2,1,107,2,5,
/* out0173_em-eta13-phi8*/	7,89,0,1,89,2,3,90,0,1,90,1,2,93,0,3,107,1,7,107,2,1,
/* out0174_em-eta14-phi8*/	4,89,0,6,93,0,2,106,2,6,107,1,1,
/* out0175_em-eta15-phi8*/	5,49,2,1,89,0,4,106,0,1,106,1,3,106,2,4,
/* out0176_em-eta16-phi8*/	3,49,1,2,49,2,3,106,1,6,
/* out0177_em-eta17-phi8*/	2,49,1,4,105,2,6,
/* out0178_em-eta18-phi8*/	3,49,1,2,105,0,4,105,2,3,
/* out0179_em-eta19-phi8*/	1,105,0,3,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	1,119,3,13,
/* out0182_em-eta2-phi9*/	2,119,2,14,119,3,3,
/* out0183_em-eta3-phi9*/	2,118,3,16,119,2,2,
/* out0184_em-eta4-phi9*/	2,94,2,2,118,2,16,
/* out0185_em-eta5-phi9*/	6,60,0,8,60,2,2,94,1,11,94,2,7,117,2,2,117,3,16,
/* out0186_em-eta6-phi9*/	7,60,0,4,93,0,2,93,1,7,93,2,14,94,1,1,116,5,2,117,2,14,
/* out0187_em-eta7-phi9*/	6,59,0,2,92,0,1,92,2,11,93,1,9,116,4,4,116,5,14,
/* out0188_em-eta8-phi9*/	5,92,0,7,92,1,9,92,2,2,116,3,4,116,4,12,
/* out0189_em-eta9-phi9*/	6,52,1,1,91,0,6,91,2,7,92,1,1,115,3,3,116,3,12,
/* out0190_em-eta10-phi9*/	5,51,2,2,91,0,9,91,1,3,115,2,3,115,3,13,
/* out0191_em-eta11-phi9*/	7,51,1,4,51,2,1,90,0,4,90,2,1,108,0,6,108,1,10,115,2,13,
/* out0192_em-eta12-phi9*/	6,50,2,2,51,1,1,90,0,6,107,0,1,107,2,9,108,1,4,
/* out0193_em-eta13-phi9*/	5,50,1,2,50,2,5,107,0,5,107,1,5,107,2,1,
/* out0194_em-eta14-phi9*/	7,50,1,6,89,0,1,90,1,1,106,0,1,106,2,3,107,0,1,107,1,3,
/* out0195_em-eta15-phi9*/	4,49,2,4,50,1,1,106,0,7,106,2,1,
/* out0196_em-eta16-phi9*/	3,49,2,4,89,2,1,106,0,5,
/* out0197_em-eta17-phi9*/	4,49,1,4,89,1,2,89,2,1,105,2,2,
/* out0198_em-eta18-phi9*/	3,49,1,3,89,1,2,105,2,3,
/* out0199_em-eta19-phi9*/	1,105,0,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	1,124,0,13,
/* out0202_em-eta2-phi10*/	2,124,0,3,124,1,14,
/* out0203_em-eta3-phi10*/	2,123,0,16,124,1,2,
/* out0204_em-eta4-phi10*/	4,55,0,1,55,1,1,94,2,3,123,1,16,
/* out0205_em-eta5-phi10*/	7,54,2,5,55,1,7,94,0,16,94,1,3,94,2,4,122,0,16,122,1,2,
/* out0206_em-eta6-phi10*/	8,53,2,1,54,1,9,54,2,3,93,0,10,93,2,2,94,1,1,121,0,2,122,1,14,
/* out0207_em-eta7-phi10*/	6,53,1,7,53,2,10,92,0,2,93,0,4,121,0,14,121,1,4,
/* out0208_em-eta8-phi10*/	5,52,2,8,53,1,5,92,0,6,121,1,12,121,2,4,
/* out0209_em-eta9-phi10*/	4,52,1,10,52,2,5,120,0,3,121,2,12,
/* out0210_em-eta10-phi10*/	5,51,2,9,52,1,3,91,0,1,120,0,13,120,1,3,
/* out0211_em-eta11-phi10*/	6,51,0,2,51,1,6,51,2,3,91,2,3,108,0,9,120,1,13,
/* out0212_em-eta12-phi10*/	6,50,2,4,51,1,5,91,1,5,91,2,4,107,0,3,108,0,1,
/* out0213_em-eta13-phi10*/	6,50,0,3,50,1,1,50,2,4,90,2,3,91,1,2,107,0,6,
/* out0214_em-eta14-phi10*/	4,50,0,2,50,1,4,90,1,3,90,2,6,
/* out0215_em-eta15-phi10*/	5,49,0,1,49,2,3,50,1,2,90,1,6,106,0,1,
/* out0216_em-eta16-phi10*/	4,49,0,3,49,2,1,89,2,6,106,0,1,
/* out0217_em-eta17-phi10*/	3,49,0,3,89,1,3,89,2,3,
/* out0218_em-eta18-phi10*/	3,49,0,2,49,1,1,89,1,5,
/* out0219_em-eta19-phi10*/	1,89,1,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	1,124,3,13,
/* out0222_em-eta2-phi11*/	2,124,2,14,124,3,3,
/* out0223_em-eta3-phi11*/	2,123,3,16,124,2,2,
/* out0224_em-eta4-phi11*/	2,55,0,2,123,2,16,
/* out0225_em-eta5-phi11*/	7,48,0,7,54,0,3,54,2,6,55,0,13,55,1,8,122,2,2,122,3,16,
/* out0226_em-eta6-phi11*/	7,47,0,4,53,2,1,54,0,13,54,1,7,54,2,2,121,5,2,122,2,14,
/* out0227_em-eta7-phi11*/	6,47,0,3,53,0,13,53,1,1,53,2,4,121,4,4,121,5,14,
/* out0228_em-eta8-phi11*/	7,46,0,6,52,0,3,52,2,3,53,0,3,53,1,3,121,3,4,121,4,12,
/* out0229_em-eta9-phi11*/	6,45,0,1,46,0,1,52,0,12,52,1,1,120,3,3,121,3,12,
/* out0230_em-eta10-phi11*/	7,45,0,6,51,0,3,51,2,1,52,0,1,52,1,1,120,2,3,120,3,13,
/* out0231_em-eta11-phi11*/	5,44,0,1,51,0,9,91,0,1,91,2,6,120,2,13,
/* out0232_em-eta12-phi11*/	7,44,0,5,50,0,1,50,2,1,51,0,2,91,0,6,91,1,4,91,2,3,
/* out0233_em-eta13-phi11*/	6,44,0,2,50,0,6,90,0,1,90,2,4,91,0,1,91,1,5,
/* out0234_em-eta14-phi11*/	5,43,0,2,50,0,4,90,0,5,90,1,1,90,2,3,
/* out0235_em-eta15-phi11*/	4,43,0,4,49,0,1,90,0,3,90,1,5,
/* out0236_em-eta16-phi11*/	4,43,0,2,49,0,3,89,0,2,89,2,4,
/* out0237_em-eta17-phi11*/	4,42,0,1,49,0,3,89,0,4,89,2,1,
/* out0238_em-eta18-phi11*/	3,42,0,3,89,0,2,89,1,2,
/* out0239_em-eta19-phi11*/	2,42,1,1,89,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	1,129,0,13,
/* out0242_em-eta2-phi12*/	2,129,0,3,129,1,14,
/* out0243_em-eta3-phi12*/	2,128,0,16,129,1,2,
/* out0244_em-eta4-phi12*/	3,41,0,1,48,1,1,128,1,16,
/* out0245_em-eta5-phi12*/	6,41,0,2,48,0,8,48,1,14,48,2,10,127,0,16,127,1,2,
/* out0246_em-eta6-phi12*/	8,40,0,1,47,0,5,47,1,14,47,2,1,48,0,1,48,2,5,126,0,2,127,1,14,
/* out0247_em-eta7-phi12*/	6,46,0,1,46,1,6,47,0,4,47,2,12,126,0,14,126,1,4,
/* out0248_em-eta8-phi12*/	5,46,0,7,46,1,6,46,2,6,126,1,12,126,2,4,
/* out0249_em-eta9-phi12*/	6,45,0,2,45,1,8,46,0,1,46,2,5,125,0,3,126,2,12,
/* out0250_em-eta10-phi12*/	5,45,0,6,45,1,2,45,2,5,125,0,13,125,1,3,
/* out0251_em-eta11-phi12*/	7,44,0,1,44,1,5,45,0,1,45,2,4,88,0,9,91,0,1,125,1,13,
/* out0252_em-eta12-phi12*/	8,44,0,5,44,1,2,44,2,1,87,0,2,87,1,1,88,0,3,88,2,2,91,0,6,
/* out0253_em-eta13-phi12*/	5,43,1,1,44,0,2,44,2,5,87,0,9,91,0,1,
/* out0254_em-eta14-phi12*/	5,43,0,2,43,1,4,87,0,3,87,2,1,90,0,5,
/* out0255_em-eta15-phi12*/	4,43,0,4,43,2,1,86,0,5,90,0,2,
/* out0256_em-eta16-phi12*/	4,43,0,2,43,2,3,86,0,5,89,0,2,
/* out0257_em-eta17-phi12*/	3,42,0,4,86,0,1,89,0,4,
/* out0258_em-eta18-phi12*/	4,42,0,3,42,1,1,85,0,3,89,0,2,
/* out0259_em-eta19-phi12*/	2,42,1,1,85,1,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	1,129,3,13,
/* out0262_em-eta2-phi13*/	2,129,2,14,129,3,3,
/* out0263_em-eta3-phi13*/	2,128,3,16,129,2,2,
/* out0264_em-eta4-phi13*/	3,41,0,5,41,2,1,128,2,16,
/* out0265_em-eta5-phi13*/	8,40,0,4,40,1,11,41,0,8,41,2,13,48,1,1,48,2,1,127,2,2,127,3,16,
/* out0266_em-eta6-phi13*/	8,39,1,3,40,0,11,40,1,1,40,2,10,47,1,2,47,2,1,126,5,2,127,2,14,
/* out0267_em-eta7-phi13*/	7,39,0,14,39,1,4,39,2,2,46,1,1,47,2,2,126,4,4,126,5,14,
/* out0268_em-eta8-phi13*/	8,38,0,4,38,1,3,39,0,2,39,2,3,46,1,3,46,2,4,126,3,4,126,4,12,
/* out0269_em-eta9-phi13*/	5,38,0,11,45,1,3,46,2,1,125,3,3,126,3,12,
/* out0270_em-eta10-phi13*/	6,37,0,3,38,2,1,45,1,3,45,2,6,125,2,3,125,3,13,
/* out0271_em-eta11-phi13*/	6,37,0,5,44,1,4,45,2,1,88,0,4,88,2,7,125,2,13,
/* out0272_em-eta12-phi13*/	5,44,1,5,44,2,4,84,0,1,87,1,8,88,2,6,
/* out0273_em-eta13-phi13*/	6,36,0,2,43,1,1,44,2,5,87,0,2,87,1,4,87,2,5,
/* out0274_em-eta14-phi13*/	3,43,1,6,86,1,3,87,2,6,
/* out0275_em-eta15-phi13*/	4,43,1,2,43,2,4,86,0,2,86,1,5,
/* out0276_em-eta16-phi13*/	3,43,2,4,86,0,3,86,2,4,
/* out0277_em-eta17-phi13*/	4,42,0,4,42,1,1,85,0,4,86,2,2,
/* out0278_em-eta18-phi13*/	4,42,0,1,42,1,3,85,0,5,85,1,2,
/* out0279_em-eta19-phi13*/	1,85,1,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	1,134,0,13,
/* out0282_em-eta2-phi14*/	2,134,0,3,134,1,14,
/* out0283_em-eta3-phi14*/	2,133,0,16,134,1,2,
/* out0284_em-eta4-phi14*/	4,24,0,4,24,2,1,41,2,1,133,1,16,
/* out0285_em-eta5-phi14*/	8,23,1,1,24,0,9,24,1,10,24,2,15,40,1,3,41,2,1,132,0,16,132,1,2,
/* out0286_em-eta6-phi14*/	8,23,0,14,23,1,4,23,2,1,39,1,2,40,1,1,40,2,6,131,0,2,132,1,14,
/* out0287_em-eta7-phi14*/	8,22,0,4,22,1,1,23,0,2,23,2,1,39,1,7,39,2,8,131,0,14,131,1,4,
/* out0288_em-eta8-phi14*/	5,22,0,5,38,1,11,39,2,3,131,1,12,131,2,4,
/* out0289_em-eta9-phi14*/	5,38,0,1,38,1,2,38,2,13,130,0,3,131,2,12,
/* out0290_em-eta10-phi14*/	5,37,0,2,37,1,10,38,2,1,130,0,13,130,1,3,
/* out0291_em-eta11-phi14*/	7,37,0,5,37,1,1,37,2,5,84,0,5,84,1,7,88,2,1,130,1,13,
/* out0292_em-eta12-phi14*/	8,36,0,2,36,1,4,37,0,1,37,2,2,44,2,1,84,0,10,84,2,2,87,1,1,
/* out0293_em-eta13-phi14*/	6,36,0,7,82,0,3,82,1,1,84,2,1,87,1,2,87,2,3,
/* out0294_em-eta14-phi14*/	5,36,0,4,43,1,1,82,0,6,86,1,2,87,2,1,
/* out0295_em-eta15-phi14*/	6,35,0,2,43,1,1,43,2,3,82,0,1,86,1,6,86,2,2,
/* out0296_em-eta16-phi14*/	3,35,0,3,43,2,1,86,2,6,
/* out0297_em-eta17-phi14*/	5,35,0,1,42,1,3,85,0,3,85,1,2,86,2,1,
/* out0298_em-eta18-phi14*/	3,42,1,4,85,0,1,85,1,5,
/* out0299_em-eta19-phi14*/	0,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	1,134,3,13,
/* out0302_em-eta2-phi15*/	2,134,2,14,134,3,3,
/* out0303_em-eta3-phi15*/	2,133,3,16,134,2,2,
/* out0304_em-eta4-phi15*/	1,133,2,16,
/* out0305_em-eta5-phi15*/	8,23,1,2,24,0,3,24,1,6,28,0,14,28,1,7,28,2,1,132,2,2,132,3,16,
/* out0306_em-eta6-phi15*/	8,23,1,9,23,2,10,26,0,4,26,1,1,28,0,2,28,2,1,131,5,2,132,2,14,
/* out0307_em-eta7-phi15*/	7,22,0,2,22,1,14,22,2,1,23,2,4,26,0,2,131,4,4,131,5,14,
/* out0308_em-eta8-phi15*/	5,21,1,2,22,0,5,22,2,10,131,3,4,131,4,12,
/* out0309_em-eta9-phi15*/	5,21,0,10,21,1,4,38,2,1,130,3,3,131,3,12,
/* out0310_em-eta10-phi15*/	6,21,0,6,21,2,1,37,1,5,37,2,1,130,2,3,130,3,13,
/* out0311_em-eta11-phi15*/	5,20,0,4,37,2,7,84,1,9,84,2,1,130,2,13,
/* out0312_em-eta12-phi15*/	5,20,0,1,36,1,7,37,2,1,83,1,1,84,2,11,
/* out0313_em-eta13-phi15*/	6,36,0,1,36,1,3,36,2,4,82,0,1,82,1,10,84,2,1,
/* out0314_em-eta14-phi15*/	5,35,1,1,36,2,6,82,0,4,82,1,1,82,2,4,
/* out0315_em-eta15-phi15*/	7,35,0,1,35,1,4,81,0,1,81,1,2,82,0,1,82,2,3,86,2,1,
/* out0316_em-eta16-phi15*/	2,35,0,4,81,0,6,
/* out0317_em-eta17-phi15*/	3,35,0,4,81,0,5,85,1,1,
/* out0318_em-eta18-phi15*/	3,35,0,1,42,1,2,85,1,4,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	1,139,0,13,
/* out0322_em-eta2-phi16*/	2,139,0,3,139,1,14,
/* out0323_em-eta3-phi16*/	2,138,0,16,139,1,2,
/* out0324_em-eta4-phi16*/	2,28,1,1,138,1,16,
/* out0325_em-eta5-phi16*/	6,27,1,7,27,2,2,28,1,8,28,2,11,137,0,16,137,1,2,
/* out0326_em-eta6-phi16*/	7,26,0,4,26,1,14,26,2,4,27,1,3,28,2,3,136,0,2,137,1,14,
/* out0327_em-eta7-phi16*/	8,22,1,1,22,2,2,25,0,2,25,1,5,26,0,6,26,2,8,136,0,14,136,1,4,
/* out0328_em-eta8-phi16*/	5,21,1,3,22,2,3,25,0,12,136,1,12,136,2,4,
/* out0329_em-eta9-phi16*/	5,21,1,7,21,2,8,25,0,1,135,0,3,136,2,12,
/* out0330_em-eta10-phi16*/	4,20,1,6,21,2,7,135,0,13,135,1,3,
/* out0331_em-eta11-phi16*/	6,20,0,6,20,1,4,20,2,1,83,1,1,83,2,6,135,1,13,
/* out0332_em-eta12-phi16*/	6,20,0,5,20,2,2,36,1,2,83,0,1,83,1,10,83,2,2,
/* out0333_em-eta13-phi16*/	6,14,1,3,36,2,4,82,1,4,82,2,1,83,0,1,83,1,4,
/* out0334_em-eta14-phi16*/	5,14,1,2,35,1,2,36,2,2,79,0,2,82,2,7,
/* out0335_em-eta15-phi16*/	4,35,1,5,79,0,1,81,1,6,82,2,1,
/* out0336_em-eta16-phi16*/	5,35,1,1,35,2,3,81,0,1,81,1,4,81,2,1,
/* out0337_em-eta17-phi16*/	3,35,2,4,81,0,2,81,2,4,
/* out0338_em-eta18-phi16*/	3,35,2,1,81,0,1,81,2,1,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	1,139,3,13,
/* out0342_em-eta2-phi17*/	2,139,2,14,139,3,3,
/* out0343_em-eta3-phi17*/	2,138,3,16,139,2,2,
/* out0344_em-eta4-phi17*/	1,138,2,16,
/* out0345_em-eta5-phi17*/	5,27,0,9,27,1,3,27,2,14,137,2,2,137,3,16,
/* out0346_em-eta6-phi17*/	8,26,1,1,26,2,2,27,0,7,27,1,3,33,0,5,33,1,8,136,5,2,137,2,14,
/* out0347_em-eta7-phi17*/	6,25,1,9,25,2,1,26,2,2,33,0,10,136,4,4,136,5,14,
/* out0348_em-eta8-phi17*/	6,25,0,1,25,1,2,25,2,14,29,2,1,136,3,4,136,4,12,
/* out0349_em-eta9-phi17*/	5,25,2,1,29,1,7,29,2,7,135,3,3,136,3,12,
/* out0350_em-eta10-phi17*/	4,20,1,3,29,1,9,135,2,3,135,3,13,
/* out0351_em-eta11-phi17*/	4,20,1,3,20,2,8,83,2,5,135,2,13,
/* out0352_em-eta12-phi17*/	4,14,2,4,20,2,5,83,0,10,83,2,3,
/* out0353_em-eta13-phi17*/	4,14,1,4,14,2,4,79,1,6,83,0,4,
/* out0354_em-eta14-phi17*/	3,14,1,6,79,0,8,79,1,1,
/* out0355_em-eta15-phi17*/	5,14,1,1,35,1,3,35,2,1,79,0,5,81,1,3,
/* out0356_em-eta16-phi17*/	3,35,2,4,81,1,1,81,2,5,
/* out0357_em-eta17-phi17*/	2,35,2,3,81,2,5,
/* out0358_em-eta18-phi17*/	0,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	1,144,0,13,
/* out0362_em-eta2-phi18*/	2,144,0,3,144,1,14,
/* out0363_em-eta3-phi18*/	2,143,0,16,144,1,2,
/* out0364_em-eta4-phi18*/	1,143,1,16,
/* out0365_em-eta5-phi18*/	5,34,0,9,34,1,14,34,2,3,142,0,16,142,1,2,
/* out0366_em-eta6-phi18*/	8,31,1,2,31,2,1,33,1,8,33,2,5,34,0,7,34,2,3,141,0,2,142,1,14,
/* out0367_em-eta7-phi18*/	7,30,1,1,30,2,9,31,1,2,33,0,1,33,2,11,141,0,14,141,1,4,
/* out0368_em-eta8-phi18*/	6,29,2,1,30,0,1,30,1,14,30,2,2,141,1,12,141,2,4,
/* out0369_em-eta9-phi18*/	5,29,0,7,29,2,7,30,1,1,140,0,3,141,2,12,
/* out0370_em-eta10-phi18*/	4,15,2,3,29,0,9,140,0,13,140,1,3,
/* out0371_em-eta11-phi18*/	4,15,1,8,15,2,3,80,1,5,140,1,13,
/* out0372_em-eta12-phi18*/	4,14,2,4,15,1,5,80,0,10,80,1,3,
/* out0373_em-eta13-phi18*/	4,14,0,4,14,2,4,79,1,7,80,0,4,
/* out0374_em-eta14-phi18*/	3,14,0,6,79,1,2,79,2,7,
/* out0375_em-eta15-phi18*/	5,7,1,1,7,2,3,14,0,1,76,2,3,79,2,5,
/* out0376_em-eta16-phi18*/	3,7,1,4,76,1,5,76,2,1,
/* out0377_em-eta17-phi18*/	2,7,1,3,76,1,5,
/* out0378_em-eta18-phi18*/	0,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	1,144,3,13,
/* out0382_em-eta2-phi19*/	2,144,2,14,144,3,3,
/* out0383_em-eta3-phi19*/	2,143,3,16,144,2,2,
/* out0384_em-eta4-phi19*/	2,32,2,1,143,2,16,
/* out0385_em-eta5-phi19*/	6,32,1,11,32,2,8,34,1,2,34,2,7,142,2,2,142,3,16,
/* out0386_em-eta6-phi19*/	7,31,0,4,31,1,4,31,2,14,32,1,3,34,2,3,141,5,2,142,2,14,
/* out0387_em-eta7-phi19*/	8,17,1,2,17,2,1,30,0,2,30,2,5,31,0,6,31,1,8,141,4,4,141,5,14,
/* out0388_em-eta8-phi19*/	5,16,2,3,17,1,3,30,0,12,141,3,4,141,4,12,
/* out0389_em-eta9-phi19*/	5,16,1,8,16,2,7,30,0,1,140,3,3,141,3,12,
/* out0390_em-eta10-phi19*/	4,15,2,6,16,1,7,140,2,3,140,3,13,
/* out0391_em-eta11-phi19*/	6,15,0,6,15,1,1,15,2,4,80,1,6,80,2,1,140,2,13,
/* out0392_em-eta12-phi19*/	6,8,2,2,15,0,5,15,1,2,80,0,1,80,1,2,80,2,10,
/* out0393_em-eta13-phi19*/	7,8,1,4,14,0,3,77,1,1,77,2,4,79,2,1,80,0,1,80,2,4,
/* out0394_em-eta14-phi19*/	5,7,2,2,8,1,2,14,0,2,77,1,7,79,2,2,
/* out0395_em-eta15-phi19*/	4,7,2,5,76,2,6,77,1,1,79,2,1,
/* out0396_em-eta16-phi19*/	5,7,1,3,7,2,1,76,0,1,76,1,1,76,2,4,
/* out0397_em-eta17-phi19*/	3,7,1,4,76,0,2,76,1,4,
/* out0398_em-eta18-phi19*/	3,7,1,1,76,0,1,76,1,1,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	1,149,0,13,
/* out0402_em-eta2-phi20*/	2,149,0,3,149,1,14,
/* out0403_em-eta3-phi20*/	2,148,0,16,149,1,2,
/* out0404_em-eta4-phi20*/	1,148,1,16,
/* out0405_em-eta5-phi20*/	8,18,2,2,19,0,3,19,2,7,32,0,14,32,1,1,32,2,7,147,0,16,147,1,2,
/* out0406_em-eta6-phi20*/	8,18,1,10,18,2,9,31,0,4,31,2,1,32,0,2,32,1,1,146,0,2,147,1,14,
/* out0407_em-eta7-phi20*/	7,17,0,2,17,1,1,17,2,14,18,1,4,31,0,2,146,0,14,146,1,4,
/* out0408_em-eta8-phi20*/	5,16,2,2,17,0,5,17,1,10,146,1,12,146,2,4,
/* out0409_em-eta9-phi20*/	5,10,1,1,16,0,10,16,2,4,145,0,3,146,2,12,
/* out0410_em-eta10-phi20*/	6,9,1,1,9,2,5,16,0,6,16,1,1,145,0,13,145,1,3,
/* out0411_em-eta11-phi20*/	5,9,1,7,15,0,4,78,1,1,78,2,9,145,1,13,
/* out0412_em-eta12-phi20*/	5,8,2,7,9,1,1,15,0,1,78,1,11,80,2,1,
/* out0413_em-eta13-phi20*/	6,8,0,1,8,1,4,8,2,3,77,0,1,77,2,10,78,1,1,
/* out0414_em-eta14-phi20*/	5,7,2,1,8,1,6,77,0,4,77,1,4,77,2,1,
/* out0415_em-eta15-phi20*/	7,7,0,1,7,2,4,73,1,1,76,0,1,76,2,2,77,0,1,77,1,3,
/* out0416_em-eta16-phi20*/	2,7,0,4,76,0,6,
/* out0417_em-eta17-phi20*/	3,7,0,4,72,1,1,76,0,5,
/* out0418_em-eta18-phi20*/	3,0,1,2,7,0,1,72,1,4,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	1,149,3,13,
/* out0422_em-eta2-phi21*/	2,149,2,14,149,3,3,
/* out0423_em-eta3-phi21*/	2,148,3,16,149,2,2,
/* out0424_em-eta4-phi21*/	4,13,1,1,19,0,4,19,1,1,148,2,16,
/* out0425_em-eta5-phi21*/	8,12,2,3,13,1,1,18,2,1,19,0,9,19,1,15,19,2,9,147,2,2,147,3,16,
/* out0426_em-eta6-phi21*/	8,11,2,2,12,1,6,12,2,1,18,0,14,18,1,1,18,2,4,146,5,2,147,2,14,
/* out0427_em-eta7-phi21*/	8,11,1,8,11,2,7,17,0,4,17,2,1,18,0,2,18,1,1,146,4,4,146,5,14,
/* out0428_em-eta8-phi21*/	5,10,2,11,11,1,3,17,0,5,146,3,4,146,4,12,
/* out0429_em-eta9-phi21*/	5,10,0,1,10,1,13,10,2,2,145,3,3,146,3,12,
/* out0430_em-eta10-phi21*/	5,9,0,2,9,2,10,10,1,1,145,2,3,145,3,13,
/* out0431_em-eta11-phi21*/	7,9,0,5,9,1,5,9,2,1,75,1,1,78,0,5,78,2,7,145,2,13,
/* out0432_em-eta12-phi21*/	8,2,1,1,8,0,2,8,2,4,9,0,1,9,1,2,74,2,1,78,0,10,78,1,2,
/* out0433_em-eta13-phi21*/	6,8,0,7,74,1,3,74,2,2,77,0,3,77,2,1,78,1,1,
/* out0434_em-eta14-phi21*/	5,1,2,1,8,0,4,73,2,2,74,1,1,77,0,6,
/* out0435_em-eta15-phi21*/	6,1,1,3,1,2,1,7,0,2,73,1,2,73,2,6,77,0,1,
/* out0436_em-eta16-phi21*/	4,0,2,1,1,1,1,7,0,3,73,1,6,
/* out0437_em-eta17-phi21*/	6,0,1,3,0,2,1,7,0,1,72,1,2,72,2,3,73,1,1,
/* out0438_em-eta18-phi21*/	3,0,1,4,72,1,5,72,2,1,
/* out0439_em-eta19-phi21*/	0,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	1,154,0,13,
/* out0442_em-eta2-phi22*/	2,154,0,3,154,1,14,
/* out0443_em-eta3-phi22*/	2,153,0,16,154,1,2,
/* out0444_em-eta4-phi22*/	3,13,0,5,13,1,1,153,1,16,
/* out0445_em-eta5-phi22*/	8,6,1,1,6,2,1,12,0,4,12,2,11,13,0,8,13,1,13,152,0,16,152,1,2,
/* out0446_em-eta6-phi22*/	8,5,1,1,5,2,2,11,2,3,12,0,11,12,1,10,12,2,1,151,0,2,152,1,14,
/* out0447_em-eta7-phi22*/	7,4,2,1,5,1,2,11,0,14,11,1,2,11,2,4,151,0,14,151,1,4,
/* out0448_em-eta8-phi22*/	8,4,1,4,4,2,3,10,0,4,10,2,3,11,0,2,11,1,3,151,1,12,151,2,4,
/* out0449_em-eta9-phi22*/	5,3,2,3,4,1,1,10,0,11,150,0,3,151,2,12,
/* out0450_em-eta10-phi22*/	6,3,1,6,3,2,3,9,0,3,10,1,1,150,0,13,150,1,3,
/* out0451_em-eta11-phi22*/	6,2,2,4,3,1,1,9,0,5,75,0,4,75,1,7,150,1,13,
/* out0452_em-eta12-phi22*/	5,2,1,4,2,2,5,74,2,8,75,1,6,78,0,1,
/* out0453_em-eta13-phi22*/	6,1,2,1,2,1,5,8,0,2,74,0,2,74,1,5,74,2,4,
/* out0454_em-eta14-phi22*/	3,1,2,6,73,2,3,74,1,6,
/* out0455_em-eta15-phi22*/	4,1,1,4,1,2,2,73,0,2,73,2,5,
/* out0456_em-eta16-phi22*/	4,0,2,1,1,1,4,73,0,3,73,1,4,
/* out0457_em-eta17-phi22*/	4,0,1,1,0,2,4,72,2,4,73,1,2,
/* out0458_em-eta18-phi22*/	4,0,1,4,0,2,1,72,1,2,72,2,5,
/* out0459_em-eta19-phi22*/	1,72,1,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	1,154,3,13,
/* out0462_em-eta2-phi23*/	2,154,2,14,154,3,3,
/* out0463_em-eta3-phi23*/	2,153,3,16,154,2,2,
/* out0464_em-eta4-phi23*/	4,6,0,7,6,2,1,13,0,1,153,2,16,
/* out0465_em-eta5-phi23*/	6,6,0,8,6,1,10,6,2,14,13,0,2,152,2,2,152,3,16,
/* out0466_em-eta6-phi23*/	8,5,0,5,5,1,1,5,2,14,6,0,1,6,1,5,12,0,1,151,5,2,152,2,14,
/* out0467_em-eta7-phi23*/	6,4,0,8,4,2,6,5,0,11,5,1,12,151,4,4,151,5,14,
/* out0468_em-eta8-phi23*/	5,4,0,7,4,1,6,4,2,6,151,3,4,151,4,12,
/* out0469_em-eta9-phi23*/	6,3,0,2,3,2,8,4,0,1,4,1,5,150,3,3,151,3,12,
/* out0470_em-eta10-phi23*/	5,3,0,13,3,1,5,3,2,2,150,2,3,150,3,13,
/* out0471_em-eta11-phi23*/	6,2,0,8,2,2,5,3,0,1,3,1,4,75,0,9,150,2,13,
/* out0472_em-eta12-phi23*/	7,2,0,6,2,1,1,2,2,2,74,0,2,74,2,1,75,0,3,75,1,2,
/* out0473_em-eta13-phi23*/	5,1,0,5,1,2,1,2,0,2,2,1,5,74,0,9,
/* out0474_em-eta14-phi23*/	4,1,0,3,1,2,4,74,0,3,74,1,1,
/* out0475_em-eta15-phi23*/	3,1,0,5,1,1,1,73,0,5,
/* out0476_em-eta16-phi23*/	3,1,0,2,1,1,3,73,0,5,
/* out0477_em-eta17-phi23*/	3,0,2,5,1,0,1,73,0,1,
/* out0478_em-eta18-phi23*/	3,0,1,1,0,2,3,72,2,3,
/* out0479_em-eta19-phi23*/	2,0,1,1,72,1,1
};