parameter integer matrixH [0:7931] = {
/* num inputs = 180(in0-in179) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 13 */
//* total number of input in adders 2483 */

/* out0000_em-eta0-phi0*/	1,135,0,10,
/* out0001_em-eta1-phi0*/	2,135,0,6,135,1,12,
/* out0002_em-eta2-phi0*/	2,134,0,14,135,1,4,
/* out0003_em-eta3-phi0*/	2,134,0,2,134,1,15,
/* out0004_em-eta4-phi0*/	2,133,0,16,134,1,1,
/* out0005_em-eta5-phi0*/	6,87,0,7,87,1,15,87,2,6,94,2,3,132,0,1,133,1,16,
/* out0006_em-eta6-phi0*/	7,86,0,10,86,1,13,87,0,9,87,2,9,93,0,1,132,0,15,132,1,3,
/* out0007_em-eta7-phi0*/	7,85,0,7,85,1,3,86,0,6,86,1,1,86,2,13,132,1,13,132,2,3,
/* out0008_em-eta8-phi0*/	5,85,0,7,85,1,9,85,2,4,269,2,5,132,2,13,
/* out0009_em-eta9-phi0*/	8,84,0,1,84,1,6,85,0,2,85,2,7,268,0,2,268,1,3,269,1,3,269,2,8,
/* out0010_em-eta10-phi0*/	5,84,0,13,84,1,4,84,2,3,268,0,12,268,1,1,
/* out0011_em-eta11-phi0*/	9,83,0,1,83,1,4,84,0,2,84,2,5,127,2,6,267,0,2,267,1,1,268,0,2,268,2,2,
/* out0012_em-eta12-phi0*/	8,83,0,6,83,1,3,83,2,1,126,0,1,126,1,1,127,1,2,127,2,6,267,0,9,
/* out0013_em-eta13-phi0*/	5,83,0,3,83,2,5,126,0,9,267,0,3,267,2,1,
/* out0014_em-eta14-phi0*/	6,82,0,2,82,1,4,83,0,6,126,0,4,126,2,1,266,0,5,
/* out0015_em-eta15-phi0*/	4,82,0,5,82,1,1,125,0,4,266,0,5,
/* out0016_em-eta16-phi0*/	5,82,0,3,82,2,2,125,0,5,265,0,1,266,0,1,
/* out0017_em-eta17-phi0*/	6,81,0,2,81,1,2,82,0,6,82,2,1,125,0,1,265,0,3,
/* out0018_em-eta18-phi0*/	3,81,0,5,124,0,3,265,0,1,
/* out0019_em-eta19-phi0*/	2,81,0,2,124,0,2,
/* out0020_em-eta0-phi1*/	1,135,3,10,
/* out0021_em-eta1-phi1*/	2,135,2,12,135,3,6,
/* out0022_em-eta2-phi1*/	2,134,3,14,135,2,4,
/* out0023_em-eta3-phi1*/	2,134,2,15,134,3,2,
/* out0024_em-eta4-phi1*/	2,133,3,16,134,2,1,
/* out0025_em-eta5-phi1*/	8,87,1,1,87,2,1,93,0,2,93,1,8,94,1,14,94,2,13,132,5,1,133,2,16,
/* out0026_em-eta6-phi1*/	6,86,1,2,93,0,13,93,1,4,93,2,10,132,4,3,132,5,15,
/* out0027_em-eta7-phi1*/	6,86,2,3,92,0,12,92,1,7,92,2,1,132,3,3,132,4,13,
/* out0028_em-eta8-phi1*/	10,85,1,4,85,2,3,91,0,2,91,1,3,92,0,4,92,2,4,263,0,1,269,1,3,269,2,3,132,3,13,
/* out0029_em-eta9-phi1*/	6,84,1,2,85,2,2,91,0,12,263,0,7,268,1,5,269,1,10,
/* out0030_em-eta10-phi1*/	7,84,1,4,84,2,5,90,0,2,91,0,1,91,2,1,268,1,7,268,2,8,
/* out0031_em-eta11-phi1*/	8,83,1,3,84,2,3,90,0,6,127,1,4,127,2,4,261,0,1,267,1,7,268,2,5,
/* out0032_em-eta12-phi1*/	9,83,1,6,83,2,3,90,0,1,122,0,1,126,1,5,127,1,9,267,0,2,267,1,5,267,2,4,
/* out0033_em-eta13-phi1*/	7,83,2,7,89,0,1,126,0,2,126,1,7,126,2,3,266,1,3,267,2,6,
/* out0034_em-eta14-phi1*/	6,82,1,6,89,0,1,125,1,2,126,2,7,266,0,2,266,1,5,
/* out0035_em-eta15-phi1*/	6,82,1,3,82,2,3,125,0,2,125,1,7,266,0,3,266,2,4,
/* out0036_em-eta16-phi1*/	6,82,2,5,125,0,3,125,2,3,265,0,1,265,1,3,266,2,3,
/* out0037_em-eta17-phi1*/	7,81,1,4,82,2,1,124,1,2,125,0,1,125,2,3,265,0,5,265,1,1,
/* out0038_em-eta18-phi1*/	5,81,0,2,81,1,3,124,0,5,124,1,1,265,0,1,
/* out0039_em-eta19-phi1*/	2,81,0,1,124,0,2,
/* out0040_em-eta0-phi2*/	1,139,0,10,
/* out0041_em-eta1-phi2*/	2,139,0,6,139,1,12,
/* out0042_em-eta2-phi2*/	2,138,0,14,139,1,4,
/* out0043_em-eta3-phi2*/	2,138,0,2,138,1,15,
/* out0044_em-eta4-phi2*/	2,137,0,16,138,1,1,
/* out0045_em-eta5-phi2*/	7,70,0,13,70,1,9,70,2,15,93,1,2,94,1,2,136,0,1,137,1,16,
/* out0046_em-eta6-phi2*/	9,69,0,12,69,1,6,70,1,1,70,2,1,92,1,1,93,1,2,93,2,6,136,0,15,136,1,3,
/* out0047_em-eta7-phi2*/	8,68,0,2,68,1,1,69,0,4,69,2,2,92,1,8,92,2,6,136,1,13,136,2,3,
/* out0048_em-eta8-phi2*/	5,68,0,6,91,1,8,92,2,5,263,1,8,136,2,13,
/* out0049_em-eta9-phi2*/	6,91,0,1,91,1,5,91,2,10,263,0,7,263,1,5,263,2,7,
/* out0050_em-eta10-phi2*/	8,90,0,1,90,1,9,91,2,4,261,0,4,261,1,7,263,0,1,263,2,3,268,2,1,
/* out0051_em-eta11-phi2*/	9,90,0,5,90,1,2,90,2,4,122,0,3,122,1,6,127,1,1,261,0,10,261,2,2,267,1,1,
/* out0052_em-eta12-phi2*/	13,89,0,1,89,1,3,90,0,1,90,2,3,122,0,11,122,1,1,122,2,2,260,0,3,260,1,1,261,0,1,261,2,1,267,1,2,267,2,3,
/* out0053_em-eta13-phi2*/	11,89,0,7,89,1,1,121,0,2,121,1,1,122,0,1,122,2,1,126,1,3,126,2,3,260,0,6,266,1,2,267,2,2,
/* out0054_em-eta14-phi2*/	8,82,1,1,89,0,5,121,0,7,125,1,1,126,2,2,260,0,1,266,1,6,266,2,1,
/* out0055_em-eta15-phi2*/	7,82,1,1,82,2,2,88,0,1,121,0,1,125,1,6,125,2,1,266,2,6,
/* out0056_em-eta16-phi2*/	5,82,2,2,88,0,3,125,2,7,265,1,5,266,2,2,
/* out0057_em-eta17-phi2*/	7,81,1,3,88,0,2,120,0,1,124,1,4,125,2,2,265,0,3,265,1,3,
/* out0058_em-eta18-phi2*/	4,81,0,2,81,1,3,124,0,2,124,1,4,
/* out0059_em-eta19-phi2*/	2,81,0,1,124,0,1,
/* out0060_em-eta0-phi3*/	1,139,3,10,
/* out0061_em-eta1-phi3*/	2,139,2,12,139,3,6,
/* out0062_em-eta2-phi3*/	2,138,3,14,139,2,4,
/* out0063_em-eta3-phi3*/	2,138,2,15,138,3,2,
/* out0064_em-eta4-phi3*/	2,137,3,16,138,2,1,
/* out0065_em-eta5-phi3*/	6,70,0,3,70,1,6,73,0,11,73,1,7,136,5,1,137,2,16,
/* out0066_em-eta6-phi3*/	8,69,1,10,69,2,8,72,0,3,72,1,1,73,0,5,73,2,2,136,4,3,136,5,15,
/* out0067_em-eta7-phi3*/	6,68,0,1,68,1,13,69,2,6,72,0,4,136,3,3,136,4,13,
/* out0068_em-eta8-phi3*/	5,68,0,7,68,1,1,68,2,11,263,1,1,136,3,13,
/* out0069_em-eta9-phi3*/	7,67,0,8,67,1,6,91,2,1,263,1,2,263,2,5,264,1,8,264,2,4,
/* out0070_em-eta10-phi3*/	7,67,0,8,67,2,1,90,1,4,261,1,9,261,2,1,263,2,1,264,1,6,
/* out0071_em-eta11-phi3*/	6,66,0,3,90,1,1,90,2,7,122,1,7,261,2,11,262,1,1,
/* out0072_em-eta12-phi3*/	9,66,0,2,89,1,6,90,2,2,122,1,2,122,2,11,123,1,1,260,0,1,260,1,10,261,2,1,
/* out0073_em-eta13-phi3*/	8,89,0,1,89,1,4,89,2,3,121,1,9,122,2,2,260,0,4,260,1,1,260,2,4,
/* out0074_em-eta14-phi3*/	8,89,2,6,121,0,4,121,1,2,121,2,3,259,0,1,259,1,2,260,0,1,260,2,3,
/* out0075_em-eta15-phi3*/	6,88,0,1,88,1,4,120,1,2,121,0,2,121,2,4,259,0,6,
/* out0076_em-eta16-phi3*/	6,88,0,4,88,1,1,120,0,5,120,1,1,259,0,5,265,1,1,
/* out0077_em-eta17-phi3*/	5,88,0,4,120,0,5,124,1,1,265,0,1,265,1,3,
/* out0078_em-eta18-phi3*/	6,81,0,1,81,1,1,88,0,1,120,0,1,124,0,1,124,1,4,
/* out0079_em-eta19-phi3*/	0,
/* out0080_em-eta0-phi4*/	1,143,0,10,
/* out0081_em-eta1-phi4*/	2,143,0,6,143,1,12,
/* out0082_em-eta2-phi4*/	2,142,0,14,143,1,4,
/* out0083_em-eta3-phi4*/	2,142,0,2,142,1,15,
/* out0084_em-eta4-phi4*/	2,141,0,16,142,1,1,
/* out0085_em-eta5-phi4*/	6,73,1,9,73,2,8,74,1,5,74,2,2,140,0,1,141,1,16,
/* out0086_em-eta6-phi4*/	7,72,0,2,72,1,14,72,2,1,73,2,6,74,1,4,140,0,15,140,1,3,
/* out0087_em-eta7-phi4*/	7,68,1,1,68,2,1,71,1,4,72,0,7,72,2,10,140,1,13,140,2,3,
/* out0088_em-eta8-phi4*/	6,67,1,1,68,2,4,71,0,12,71,1,2,264,2,1,140,2,13,
/* out0089_em-eta9-phi4*/	6,67,1,9,67,2,6,71,0,2,264,0,6,264,1,1,264,2,11,
/* out0090_em-eta10-phi4*/	5,66,1,4,67,2,9,262,2,5,264,0,9,264,1,1,
/* out0091_em-eta11-phi4*/	6,66,0,5,66,1,6,66,2,1,123,2,4,262,1,10,262,2,3,
/* out0092_em-eta12-phi4*/	10,66,0,6,66,2,2,89,1,1,123,0,1,123,1,9,123,2,4,260,1,4,260,2,1,262,0,1,262,1,5,
/* out0093_em-eta13-phi4*/	8,60,1,2,89,1,1,89,2,4,121,1,4,123,0,1,123,1,6,260,2,7,270,1,2,
/* out0094_em-eta14-phi4*/	8,60,1,2,88,1,1,89,2,3,116,0,2,121,2,7,259,1,6,260,2,1,270,1,1,
/* out0095_em-eta15-phi4*/	7,88,1,5,116,0,1,120,1,5,121,2,2,259,0,1,259,1,4,259,2,1,
/* out0096_em-eta16-phi4*/	7,88,1,2,88,2,2,120,0,1,120,1,5,120,2,1,259,0,2,259,2,4,
/* out0097_em-eta17-phi4*/	5,88,2,4,120,0,2,120,2,3,259,0,1,259,2,1,
/* out0098_em-eta18-phi4*/	3,88,2,2,120,0,1,120,2,2,
/* out0099_em-eta19-phi4*/	0,
/* out0100_em-eta0-phi5*/	1,143,3,10,
/* out0101_em-eta1-phi5*/	2,143,2,12,143,3,6,
/* out0102_em-eta2-phi5*/	2,142,3,14,143,2,4,
/* out0103_em-eta3-phi5*/	2,142,2,15,142,3,2,
/* out0104_em-eta4-phi5*/	2,141,3,16,142,2,1,
/* out0105_em-eta5-phi5*/	5,74,0,6,74,1,2,74,2,14,140,5,1,141,2,16,
/* out0106_em-eta6-phi5*/	8,72,1,1,72,2,2,74,0,10,74,1,5,77,0,3,77,1,8,140,4,3,140,5,15,
/* out0107_em-eta7-phi5*/	5,71,1,6,72,2,3,77,0,13,140,3,3,140,4,13,
/* out0108_em-eta8-phi5*/	4,71,0,1,71,1,4,71,2,13,140,3,13,
/* out0109_em-eta9-phi5*/	7,71,0,1,71,2,3,75,1,4,75,2,8,264,0,1,272,0,6,272,1,8,
/* out0110_em-eta10-phi5*/	4,66,1,2,75,1,11,262,2,5,272,0,10,
/* out0111_em-eta11-phi5*/	5,66,1,4,66,2,6,123,2,3,262,0,10,262,2,3,
/* out0112_em-eta12-phi5*/	6,60,2,2,66,2,7,123,0,8,123,2,5,262,0,5,270,2,6,
/* out0113_em-eta13-phi5*/	6,60,1,3,60,2,5,116,1,5,123,0,6,270,1,8,270,2,2,
/* out0114_em-eta14-phi5*/	5,60,1,7,116,0,7,116,1,3,259,1,2,270,1,5,
/* out0115_em-eta15-phi5*/	7,60,1,2,88,1,3,88,2,1,116,0,6,120,1,1,259,1,2,259,2,5,
/* out0116_em-eta16-phi5*/	4,88,2,4,120,1,2,120,2,4,259,2,5,
/* out0117_em-eta17-phi5*/	2,88,2,3,120,2,5,
/* out0118_em-eta18-phi5*/	1,120,2,1,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	1,147,0,10,
/* out0121_em-eta1-phi6*/	2,147,0,6,147,1,12,
/* out0122_em-eta2-phi6*/	2,146,0,14,147,1,4,
/* out0123_em-eta3-phi6*/	2,146,0,2,146,1,15,
/* out0124_em-eta4-phi6*/	2,145,0,16,146,1,1,
/* out0125_em-eta5-phi6*/	5,79,0,6,79,1,14,79,2,2,144,0,1,145,1,16,
/* out0126_em-eta6-phi6*/	8,77,1,8,77,2,3,78,1,2,78,2,1,79,0,10,79,2,5,144,0,15,144,1,3,
/* out0127_em-eta7-phi6*/	5,76,2,6,77,2,13,78,1,3,144,1,13,144,2,3,
/* out0128_em-eta8-phi6*/	4,76,0,1,76,1,13,76,2,4,144,2,13,
/* out0129_em-eta9-phi6*/	7,75,0,5,75,2,8,76,0,1,76,1,3,272,1,8,272,2,5,273,1,1,
/* out0130_em-eta10-phi6*/	5,61,2,2,75,0,11,75,1,1,271,2,5,272,2,11,
/* out0131_em-eta11-phi6*/	5,61,1,6,61,2,4,118,1,3,271,1,10,271,2,3,
/* out0132_em-eta12-phi6*/	6,60,2,2,61,1,7,118,0,8,118,1,5,270,2,6,271,1,5,
/* out0133_em-eta13-phi6*/	6,60,0,3,60,2,6,116,1,5,118,0,6,270,0,7,270,2,2,
/* out0134_em-eta14-phi6*/	5,60,0,6,116,1,3,116,2,6,255,2,2,270,0,5,
/* out0135_em-eta15-phi6*/	7,53,1,1,53,2,3,60,0,2,115,2,1,116,2,6,255,1,5,255,2,2,
/* out0136_em-eta16-phi6*/	4,53,1,4,115,1,4,115,2,2,255,1,5,
/* out0137_em-eta17-phi6*/	2,53,1,3,115,1,5,
/* out0138_em-eta18-phi6*/	1,115,1,1,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	1,147,3,10,
/* out0141_em-eta1-phi7*/	2,147,2,12,147,3,6,
/* out0142_em-eta2-phi7*/	2,146,3,14,147,2,4,
/* out0143_em-eta3-phi7*/	2,146,2,15,146,3,2,
/* out0144_em-eta4-phi7*/	2,145,3,16,146,2,1,
/* out0145_em-eta5-phi7*/	6,79,1,2,79,2,5,80,1,8,80,2,9,144,5,1,145,2,16,
/* out0146_em-eta6-phi7*/	7,78,0,2,78,1,1,78,2,14,79,2,4,80,1,6,144,4,3,144,5,15,
/* out0147_em-eta7-phi7*/	7,63,1,1,63,2,1,76,2,4,78,0,7,78,1,10,144,3,3,144,4,13,
/* out0148_em-eta8-phi7*/	6,62,2,1,63,1,4,76,0,12,76,2,2,273,2,1,144,3,13,
/* out0149_em-eta9-phi7*/	6,62,1,6,62,2,9,76,0,2,273,0,1,273,1,6,273,2,11,
/* out0150_em-eta10-phi7*/	6,61,2,4,62,1,9,271,0,1,271,2,5,273,0,1,273,1,9,
/* out0151_em-eta11-phi7*/	6,61,0,5,61,1,1,61,2,6,118,1,4,271,0,10,271,2,3,
/* out0152_em-eta12-phi7*/	10,54,2,1,61,0,6,61,1,2,118,0,1,118,1,4,118,2,9,256,1,1,256,2,4,271,0,4,271,1,1,
/* out0153_em-eta13-phi7*/	9,54,1,4,54,2,1,60,0,2,60,2,1,117,2,4,118,0,1,118,2,6,256,1,7,270,0,3,
/* out0154_em-eta14-phi7*/	8,53,2,1,54,1,3,60,0,3,116,2,3,117,1,7,255,2,6,256,1,1,270,0,1,
/* out0155_em-eta15-phi7*/	7,53,2,5,115,2,5,116,2,1,117,1,2,255,0,1,255,1,1,255,2,4,
/* out0156_em-eta16-phi7*/	7,53,1,2,53,2,2,115,0,1,115,1,1,115,2,5,255,0,2,255,1,4,
/* out0157_em-eta17-phi7*/	5,53,1,4,115,0,2,115,1,3,255,0,1,255,1,1,
/* out0158_em-eta18-phi7*/	3,53,1,2,115,0,1,115,1,2,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	1,151,0,10,
/* out0161_em-eta1-phi8*/	2,151,0,6,151,1,12,
/* out0162_em-eta2-phi8*/	2,150,0,14,151,1,4,
/* out0163_em-eta3-phi8*/	2,150,0,2,150,1,15,
/* out0164_em-eta4-phi8*/	2,149,0,16,150,1,1,
/* out0165_em-eta5-phi8*/	6,65,0,3,65,2,7,80,0,11,80,2,7,148,0,1,149,1,16,
/* out0166_em-eta6-phi8*/	8,64,1,8,64,2,10,78,0,3,78,2,1,80,0,5,80,1,2,148,0,15,148,1,3,
/* out0167_em-eta7-phi8*/	6,63,0,1,63,2,13,64,1,6,78,0,4,148,1,13,148,2,3,
/* out0168_em-eta8-phi8*/	5,63,0,7,63,1,11,63,2,1,258,2,1,148,2,13,
/* out0169_em-eta9-phi8*/	7,56,1,1,62,0,8,62,2,6,258,1,5,258,2,2,273,0,8,273,2,4,
/* out0170_em-eta10-phi8*/	7,55,2,4,62,0,8,62,1,1,257,1,1,257,2,9,258,1,1,273,0,6,
/* out0171_em-eta11-phi8*/	6,55,1,7,55,2,1,61,0,3,119,2,7,257,1,11,271,0,1,
/* out0172_em-eta12-phi8*/	9,54,2,6,55,1,2,61,0,2,118,2,1,119,1,11,119,2,2,256,0,1,256,2,10,257,1,1,
/* out0173_em-eta13-phi8*/	8,54,0,1,54,1,3,54,2,4,117,2,9,119,1,2,256,0,4,256,1,4,256,2,1,
/* out0174_em-eta14-phi8*/	8,54,1,6,117,0,4,117,1,3,117,2,2,255,0,1,255,2,2,256,0,1,256,1,3,
/* out0175_em-eta15-phi8*/	6,53,0,1,53,2,4,115,2,2,117,0,2,117,1,4,255,0,6,
/* out0176_em-eta16-phi8*/	6,53,0,4,53,2,1,115,0,5,115,2,1,250,1,1,255,0,5,
/* out0177_em-eta17-phi8*/	3,53,0,4,115,0,5,250,1,4,
/* out0178_em-eta18-phi8*/	4,46,1,2,53,0,1,111,1,5,115,0,1,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	1,151,3,10,
/* out0181_em-eta1-phi9*/	2,151,2,12,151,3,6,
/* out0182_em-eta2-phi9*/	2,150,3,14,151,2,4,
/* out0183_em-eta3-phi9*/	2,150,2,15,150,3,2,
/* out0184_em-eta4-phi9*/	2,149,3,16,150,2,1,
/* out0185_em-eta5-phi9*/	7,58,2,2,59,1,2,65,0,13,65,1,15,65,2,7,148,5,1,149,2,16,
/* out0186_em-eta6-phi9*/	9,57,2,1,58,1,6,58,2,2,64,0,12,64,2,6,65,1,1,65,2,2,148,4,3,148,5,15,
/* out0187_em-eta7-phi9*/	8,57,1,6,57,2,8,63,0,2,63,2,1,64,0,4,64,1,2,148,3,3,148,4,13,
/* out0188_em-eta8-phi9*/	5,56,2,8,57,1,5,63,0,6,258,2,8,148,3,13,
/* out0189_em-eta9-phi9*/	6,56,0,1,56,1,10,56,2,5,258,0,7,258,1,7,258,2,5,
/* out0190_em-eta10-phi9*/	8,55,0,1,55,2,9,56,1,4,253,1,1,257,0,4,257,2,7,258,0,1,258,1,3,
/* out0191_em-eta11-phi9*/	9,55,0,5,55,1,4,55,2,2,114,1,1,119,0,3,119,2,6,252,2,1,257,0,10,257,1,2,
/* out0192_em-eta12-phi9*/	13,54,0,1,54,2,3,55,0,1,55,1,3,119,0,11,119,1,2,119,2,1,252,1,3,252,2,2,256,0,3,256,2,1,257,0,1,257,1,1,
/* out0193_em-eta13-phi9*/	11,54,0,7,54,2,1,113,1,3,113,2,3,117,0,2,117,2,1,119,0,1,119,1,1,251,2,2,252,1,2,256,0,6,
/* out0194_em-eta14-phi9*/	8,47,2,1,54,0,5,112,2,1,113,1,2,117,0,7,251,1,1,251,2,6,256,0,1,
/* out0195_em-eta15-phi9*/	7,47,1,2,47,2,1,53,0,1,112,1,1,112,2,6,117,0,1,251,1,6,
/* out0196_em-eta16-phi9*/	6,47,1,2,53,0,3,112,1,7,250,1,2,250,2,2,251,1,2,
/* out0197_em-eta17-phi9*/	8,46,1,2,53,0,2,111,1,1,111,2,2,112,1,2,115,0,1,250,1,5,250,2,1,
/* out0198_em-eta18-phi9*/	4,46,1,4,111,1,5,111,2,1,250,1,1,
/* out0199_em-eta19-phi9*/	1,111,1,1,
/* out0200_em-eta0-phi10*/	1,155,0,10,
/* out0201_em-eta1-phi10*/	2,155,0,6,155,1,12,
/* out0202_em-eta2-phi10*/	2,154,0,14,155,1,4,
/* out0203_em-eta3-phi10*/	2,154,0,2,154,1,15,
/* out0204_em-eta4-phi10*/	2,153,0,16,154,1,1,
/* out0205_em-eta5-phi10*/	8,52,1,1,52,2,1,58,0,2,58,2,8,59,0,13,59,1,14,152,0,1,153,1,16,
/* out0206_em-eta6-phi10*/	6,51,2,2,58,0,13,58,1,10,58,2,4,152,0,15,152,1,3,
/* out0207_em-eta7-phi10*/	6,51,1,3,57,0,12,57,1,1,57,2,7,152,1,13,152,2,3,
/* out0208_em-eta8-phi10*/	10,50,1,3,50,2,4,56,0,2,56,2,3,57,0,4,57,1,4,254,0,3,254,1,3,258,0,1,152,2,13,
/* out0209_em-eta9-phi10*/	6,49,2,2,50,1,2,56,0,12,253,2,5,254,1,10,258,0,7,
/* out0210_em-eta10-phi10*/	7,49,1,5,49,2,4,55,0,2,56,0,1,56,1,1,253,1,8,253,2,7,
/* out0211_em-eta11-phi10*/	8,48,2,3,49,1,3,55,0,6,114,0,4,114,1,4,252,2,7,253,1,5,257,0,1,
/* out0212_em-eta12-phi10*/	9,48,1,3,48,2,6,55,0,1,113,2,5,114,1,9,119,0,1,252,0,2,252,1,4,252,2,5,
/* out0213_em-eta13-phi10*/	7,48,1,7,54,0,1,113,0,2,113,1,3,113,2,7,251,2,3,252,1,6,
/* out0214_em-eta14-phi10*/	6,47,2,6,54,0,1,112,2,2,113,1,7,251,0,2,251,2,5,
/* out0215_em-eta15-phi10*/	6,47,1,3,47,2,3,112,0,2,112,2,7,251,0,3,251,1,4,
/* out0216_em-eta16-phi10*/	5,47,1,5,112,0,3,112,1,3,250,2,4,251,1,3,
/* out0217_em-eta17-phi10*/	8,46,1,1,46,2,3,47,1,1,111,2,3,112,0,1,112,1,3,250,1,1,250,2,5,
/* out0218_em-eta18-phi10*/	5,46,1,3,46,2,1,111,1,1,111,2,6,250,1,1,
/* out0219_em-eta19-phi10*/	2,46,1,1,111,1,2,
/* out0220_em-eta0-phi11*/	1,155,3,10,
/* out0221_em-eta1-phi11*/	2,155,2,12,155,3,6,
/* out0222_em-eta2-phi11*/	2,154,3,14,155,2,4,
/* out0223_em-eta3-phi11*/	2,154,2,15,154,3,2,
/* out0224_em-eta4-phi11*/	2,153,3,16,154,2,1,
/* out0225_em-eta5-phi11*/	6,52,0,7,52,1,6,52,2,15,59,0,3,152,5,1,153,2,16,
/* out0226_em-eta6-phi11*/	7,51,0,3,51,2,13,52,0,2,52,1,9,58,0,1,152,4,3,152,5,15,
/* out0227_em-eta7-phi11*/	6,50,2,3,51,0,5,51,1,13,51,2,1,152,3,3,152,4,13,
/* out0228_em-eta8-phi11*/	5,50,0,7,50,1,4,50,2,9,254,0,5,152,3,13,
/* out0229_em-eta9-phi11*/	9,49,0,1,49,2,6,50,0,2,50,1,7,249,0,6,253,0,2,253,2,3,254,0,8,254,1,3,
/* out0230_em-eta10-phi11*/	7,49,0,6,49,1,3,49,2,4,248,0,1,249,0,1,253,0,12,253,2,1,
/* out0231_em-eta11-phi11*/	10,48,0,1,48,2,4,49,0,1,49,1,5,114,0,6,248,0,6,252,0,2,252,2,1,253,0,2,253,1,2,
/* out0232_em-eta12-phi11*/	10,48,0,5,48,1,1,48,2,3,110,0,6,113,0,1,113,2,1,114,0,6,114,1,2,248,0,1,252,0,9,
/* out0233_em-eta13-phi11*/	7,48,0,3,48,1,5,110,0,2,113,0,9,247,0,5,252,0,3,252,1,1,
/* out0234_em-eta14-phi11*/	7,47,0,2,47,2,4,109,0,4,113,0,4,113,1,1,247,0,2,251,0,5,
/* out0235_em-eta15-phi11*/	6,47,0,4,47,2,1,109,0,3,112,0,4,246,0,2,251,0,5,
/* out0236_em-eta16-phi11*/	6,47,0,2,47,1,2,108,0,1,112,0,5,246,0,4,251,0,1,
/* out0237_em-eta17-phi11*/	6,46,2,4,47,1,1,108,0,4,112,0,1,246,0,2,250,2,3,
/* out0238_em-eta18-phi11*/	6,46,1,1,46,2,4,108,0,3,111,2,3,250,1,1,250,2,1,
/* out0239_em-eta19-phi11*/	3,46,1,1,111,1,1,111,2,1,
/* out0240_em-eta0-phi12*/	1,159,0,10,
/* out0241_em-eta1-phi12*/	2,159,0,6,159,1,12,
/* out0242_em-eta2-phi12*/	2,158,0,14,159,1,4,
/* out0243_em-eta3-phi12*/	2,158,0,2,158,1,15,
/* out0244_em-eta4-phi12*/	2,157,0,16,158,1,1,
/* out0245_em-eta5-phi12*/	7,44,0,1,44,1,5,45,0,14,45,2,8,52,0,6,156,0,1,157,1,16,
/* out0246_em-eta6-phi12*/	7,44,0,15,44,1,3,44,2,6,51,0,3,52,0,1,156,0,15,156,1,3,
/* out0247_em-eta7-phi12*/	6,43,0,11,43,1,5,44,2,1,51,0,5,156,1,13,156,2,3,
/* out0248_em-eta8-phi12*/	7,42,0,1,42,1,2,43,0,5,43,2,4,50,0,6,249,1,3,156,2,13,
/* out0249_em-eta9-phi12*/	7,42,0,12,42,1,1,49,0,1,50,0,1,249,0,7,249,1,9,249,2,4,
/* out0250_em-eta10-phi12*/	9,41,0,2,41,1,1,42,0,2,42,2,2,49,0,6,248,0,1,248,1,6,249,0,2,249,2,7,
/* out0251_em-eta11-phi12*/	6,41,0,9,49,0,1,110,1,5,248,0,6,248,1,4,248,2,3,
/* out0252_em-eta12-phi12*/	10,41,0,3,41,2,1,48,0,5,110,0,6,110,1,5,110,2,2,247,0,1,247,1,4,248,0,1,248,2,5,
/* out0253_em-eta13-phi12*/	8,40,0,5,48,0,2,109,1,3,110,0,2,110,2,6,247,0,5,247,1,3,247,2,1,
/* out0254_em-eta14-phi12*/	6,40,0,5,47,0,2,109,0,5,109,1,4,247,0,3,247,2,5,
/* out0255_em-eta15-phi12*/	7,40,0,1,47,0,4,109,0,4,109,2,5,246,0,2,246,1,4,247,2,1,
/* out0256_em-eta16-phi12*/	7,39,0,3,47,0,2,108,0,1,108,1,4,109,2,1,246,0,4,246,1,1,
/* out0257_em-eta17-phi12*/	6,39,0,3,46,2,1,108,0,4,108,1,1,246,0,2,246,2,2,
/* out0258_em-eta18-phi12*/	5,39,0,1,46,2,3,108,0,3,108,2,2,246,2,1,
/* out0259_em-eta19-phi12*/	2,46,1,1,108,2,2,
/* out0260_em-eta0-phi13*/	1,159,3,10,
/* out0261_em-eta1-phi13*/	2,159,2,12,159,3,6,
/* out0262_em-eta2-phi13*/	2,158,3,14,159,2,4,
/* out0263_em-eta3-phi13*/	2,158,2,15,158,3,2,
/* out0264_em-eta4-phi13*/	2,157,3,16,158,2,1,
/* out0265_em-eta5-phi13*/	8,38,0,14,38,1,7,38,2,2,44,1,3,45,0,2,45,2,8,156,5,1,157,2,16,
/* out0266_em-eta6-phi13*/	8,37,0,7,37,1,2,38,0,2,38,2,2,44,1,5,44,2,9,156,4,3,156,5,15,
/* out0267_em-eta7-phi13*/	6,36,0,1,37,0,7,43,1,11,43,2,4,156,3,3,156,4,13,
/* out0268_em-eta8-phi13*/	5,36,0,7,42,1,5,43,2,8,245,0,7,156,3,13,
/* out0269_em-eta9-phi13*/	9,42,0,1,42,1,8,42,2,8,244,0,2,244,1,3,245,0,6,245,2,4,249,1,4,249,2,3,
/* out0270_em-eta10-phi13*/	6,35,0,1,41,1,7,42,2,5,244,0,12,248,1,2,249,2,2,
/* out0271_em-eta11-phi13*/	10,41,0,2,41,1,5,41,2,4,107,0,7,110,1,1,243,0,2,244,0,1,244,2,1,248,1,4,248,2,5,
/* out0272_em-eta12-phi13*/	9,40,1,3,41,2,6,105,0,2,107,0,4,110,1,5,110,2,4,243,0,6,247,1,3,248,2,3,
/* out0273_em-eta13-phi13*/	8,40,0,2,40,1,5,105,0,6,109,1,2,110,2,4,243,0,1,247,1,6,247,2,3,
/* out0274_em-eta14-phi13*/	7,40,0,3,40,2,4,105,0,1,109,1,7,109,2,2,242,0,1,247,2,6,
/* out0275_em-eta15-phi13*/	6,39,1,2,40,2,3,103,0,1,109,2,7,242,0,1,246,1,6,
/* out0276_em-eta16-phi13*/	7,39,0,3,39,1,2,103,0,1,108,1,5,109,2,1,246,1,3,246,2,3,
/* out0277_em-eta17-phi13*/	4,39,0,4,108,1,4,108,2,2,246,2,5,
/* out0278_em-eta18-phi13*/	4,39,0,2,39,2,1,108,2,5,246,2,1,
/* out0279_em-eta19-phi13*/	2,39,2,1,108,2,1,
/* out0280_em-eta0-phi14*/	1,163,0,10,
/* out0281_em-eta1-phi14*/	2,163,0,6,163,1,12,
/* out0282_em-eta2-phi14*/	2,162,0,14,163,1,4,
/* out0283_em-eta3-phi14*/	2,162,0,2,162,1,15,
/* out0284_em-eta4-phi14*/	2,161,0,16,162,1,1,
/* out0285_em-eta5-phi14*/	6,32,0,6,32,1,2,38,1,9,38,2,9,160,0,1,161,1,16,
/* out0286_em-eta6-phi14*/	7,32,0,7,37,0,1,37,1,14,37,2,4,38,2,3,160,0,15,160,1,3,
/* out0287_em-eta7-phi14*/	6,31,0,3,36,1,8,37,0,1,37,2,12,160,1,13,160,2,3,
/* out0288_em-eta8-phi14*/	8,36,0,7,36,1,5,36,2,7,240,0,1,240,2,3,245,0,3,245,2,5,160,2,13,
/* out0289_em-eta9-phi14*/	8,35,0,4,35,1,6,36,0,1,36,2,3,42,2,1,240,2,7,244,1,8,245,2,7,
/* out0290_em-eta10-phi14*/	6,35,0,10,35,2,2,41,1,1,244,0,1,244,1,4,244,2,11,
/* out0291_em-eta11-phi14*/	11,34,0,3,34,1,1,35,0,1,35,2,1,41,1,2,41,2,3,107,0,5,107,2,7,243,0,1,243,1,9,244,2,3,
/* out0292_em-eta12-phi14*/	8,34,0,6,40,1,2,41,2,2,105,1,8,107,2,7,243,0,5,243,1,2,243,2,4,
/* out0293_em-eta13-phi14*/	10,34,0,1,40,1,6,40,2,1,105,0,5,105,1,3,105,2,3,242,0,1,242,1,3,243,0,1,243,2,3,
/* out0294_em-eta14-phi14*/	6,40,2,6,103,1,3,105,0,2,105,2,4,242,0,7,242,1,1,
/* out0295_em-eta15-phi14*/	6,39,1,4,40,2,2,103,0,7,103,1,1,242,0,5,246,1,1,
/* out0296_em-eta16-phi14*/	5,39,1,4,103,0,6,241,1,1,246,1,1,246,2,2,
/* out0297_em-eta17-phi14*/	8,39,2,4,102,1,1,103,0,1,103,2,1,108,1,2,108,2,2,241,1,3,246,2,2,
/* out0298_em-eta18-phi14*/	4,39,2,3,102,1,2,108,2,2,241,0,1,
/* out0299_em-eta19-phi14*/	2,102,0,1,102,1,1,
/* out0300_em-eta0-phi15*/	1,163,3,10,
/* out0301_em-eta1-phi15*/	2,163,2,12,163,3,6,
/* out0302_em-eta2-phi15*/	2,162,3,14,163,2,4,
/* out0303_em-eta3-phi15*/	2,162,2,15,162,3,2,
/* out0304_em-eta4-phi15*/	3,28,0,1,161,3,16,162,2,1,
/* out0305_em-eta5-phi15*/	9,26,0,1,28,0,10,28,1,1,28,2,16,32,0,1,32,1,14,32,2,3,160,5,1,161,2,16,
/* out0306_em-eta6-phi15*/	7,26,0,2,31,0,1,31,1,10,32,0,2,32,2,13,160,4,3,160,5,15,
/* out0307_em-eta7-phi15*/	6,31,0,12,31,1,3,31,2,7,36,1,1,160,3,3,160,4,13,
/* out0308_em-eta8-phi15*/	7,30,0,8,30,1,4,31,2,1,36,1,2,36,2,5,240,0,11,160,3,13,
/* out0309_em-eta9-phi15*/	7,30,0,6,35,1,9,35,2,1,36,2,1,240,0,3,240,1,11,240,2,6,
/* out0310_em-eta10-phi15*/	7,29,0,1,35,1,1,35,2,11,238,0,8,238,1,6,244,1,1,244,2,1,
/* out0311_em-eta11-phi15*/	9,34,0,1,34,1,10,35,2,1,106,0,8,106,2,6,107,2,2,238,0,8,238,2,1,243,1,4,
/* out0312_em-eta12-phi15*/	9,34,0,4,34,1,1,34,2,4,105,1,3,106,1,2,106,2,10,237,0,3,243,1,1,243,2,7,
/* out0313_em-eta13-phi15*/	10,33,0,1,33,1,2,34,0,1,34,2,3,104,1,3,105,1,2,105,2,6,237,0,2,242,1,6,243,2,2,
/* out0314_em-eta14-phi15*/	7,33,0,6,103,1,5,104,1,2,105,2,3,242,0,1,242,1,4,242,2,3,
/* out0315_em-eta15-phi15*/	5,33,0,5,39,1,1,103,1,5,103,2,2,242,2,6,
/* out0316_em-eta16-phi15*/	4,39,1,3,39,2,1,103,2,6,241,1,5,
/* out0317_em-eta17-phi15*/	5,39,2,4,102,1,4,103,2,1,241,0,2,241,1,3,
/* out0318_em-eta18-phi15*/	4,39,2,2,102,0,1,102,1,4,241,0,3,
/* out0319_em-eta19-phi15*/	1,102,0,4,
/* out0320_em-eta0-phi16*/	1,167,0,10,
/* out0321_em-eta1-phi16*/	2,167,0,6,167,1,12,
/* out0322_em-eta2-phi16*/	2,166,0,14,167,1,4,
/* out0323_em-eta3-phi16*/	2,166,0,2,166,1,15,
/* out0324_em-eta4-phi16*/	2,165,0,16,166,1,1,
/* out0325_em-eta5-phi16*/	9,26,0,1,26,1,12,27,0,2,27,1,13,27,2,1,28,0,5,28,1,15,164,0,1,165,1,16,
/* out0326_em-eta6-phi16*/	7,25,1,1,26,0,12,26,1,2,26,2,10,31,1,2,164,0,15,164,1,3,
/* out0327_em-eta7-phi16*/	7,25,0,11,25,1,3,30,1,1,31,1,1,31,2,8,164,1,13,164,2,3,
/* out0328_em-eta8-phi16*/	8,25,0,2,30,0,1,30,1,11,30,2,5,239,0,3,240,0,1,240,1,1,164,2,13,
/* out0329_em-eta9-phi16*/	7,29,1,5,30,0,1,30,2,9,238,1,1,239,0,4,239,2,14,240,1,4,
/* out0330_em-eta10-phi16*/	5,29,0,10,29,1,3,238,1,9,238,2,6,239,2,2,
/* out0331_em-eta11-phi16*/	8,29,0,5,29,2,1,34,1,4,34,2,1,106,0,8,106,1,4,237,1,4,238,2,9,
/* out0332_em-eta12-phi16*/	7,14,1,2,34,2,7,104,2,2,106,1,10,237,0,5,237,1,6,237,2,1,
/* out0333_em-eta13-phi16*/	8,14,1,1,33,1,6,34,2,1,104,1,4,104,2,7,237,0,6,237,2,2,242,1,1,
/* out0334_em-eta14-phi16*/	8,33,0,1,33,1,4,33,2,1,104,0,2,104,1,7,231,1,2,242,1,1,242,2,4,
/* out0335_em-eta15-phi16*/	9,33,0,2,33,2,4,98,1,1,103,1,2,103,2,3,104,0,1,231,1,2,241,1,1,242,2,3,
/* out0336_em-eta16-phi16*/	7,0,1,2,33,0,1,33,2,1,98,1,3,103,2,3,241,1,2,241,2,3,
/* out0337_em-eta17-phi16*/	6,0,1,3,102,1,2,102,2,3,241,0,3,241,1,1,241,2,2,
/* out0338_em-eta18-phi16*/	6,0,0,2,0,1,2,102,0,2,102,1,2,102,2,2,241,0,4,
/* out0339_em-eta19-phi16*/	1,102,0,6,
/* out0340_em-eta0-phi17*/	1,167,3,10,
/* out0341_em-eta1-phi17*/	2,167,2,12,167,3,6,
/* out0342_em-eta2-phi17*/	2,166,3,14,167,2,4,
/* out0343_em-eta3-phi17*/	2,166,2,15,166,3,2,
/* out0344_em-eta4-phi17*/	2,165,3,16,166,2,1,
/* out0345_em-eta5-phi17*/	7,23,1,5,26,1,2,27,0,14,27,1,3,27,2,15,164,5,1,165,2,16,
/* out0346_em-eta6-phi17*/	6,23,0,15,23,1,2,25,1,4,26,2,6,164,4,3,164,5,15,
/* out0347_em-eta7-phi17*/	5,25,0,2,25,1,8,25,2,13,164,3,3,164,4,13,
/* out0348_em-eta8-phi17*/	7,19,1,5,19,2,8,25,0,1,25,2,3,30,2,1,239,0,2,164,3,13,
/* out0349_em-eta9-phi17*/	5,19,1,11,29,1,5,30,2,1,239,0,7,239,1,13,
/* out0350_em-eta10-phi17*/	5,29,1,3,29,2,10,235,0,5,235,1,8,239,1,3,
/* out0351_em-eta11-phi17*/	6,14,2,6,29,2,5,101,0,8,101,2,2,235,0,11,237,1,2,
/* out0352_em-eta12-phi17*/	8,14,1,8,14,2,2,101,0,1,101,1,1,101,2,13,104,2,1,237,1,4,237,2,6,
/* out0353_em-eta13-phi17*/	7,14,1,5,33,1,2,101,2,1,104,0,5,104,2,6,231,2,2,237,2,7,
/* out0354_em-eta14-phi17*/	6,33,1,2,33,2,5,98,2,1,104,0,8,231,1,3,231,2,5,
/* out0355_em-eta15-phi17*/	4,33,2,5,98,1,2,98,2,6,231,1,7,
/* out0356_em-eta16-phi17*/	4,0,1,4,98,1,7,231,1,2,241,2,4,
/* out0357_em-eta17-phi17*/	4,0,1,3,98,1,3,102,2,3,241,2,5,
/* out0358_em-eta18-phi17*/	4,0,0,4,102,2,6,241,0,3,241,2,2,
/* out0359_em-eta19-phi17*/	2,102,0,2,102,2,2,
/* out0360_em-eta0-phi18*/	1,171,0,10,
/* out0361_em-eta1-phi18*/	2,171,0,6,171,1,12,
/* out0362_em-eta2-phi18*/	2,170,0,14,171,1,4,
/* out0363_em-eta3-phi18*/	2,170,0,2,170,1,15,
/* out0364_em-eta4-phi18*/	2,169,0,16,170,1,1,
/* out0365_em-eta5-phi18*/	7,21,2,2,23,1,6,24,0,15,24,1,9,24,2,16,168,0,1,169,1,16,
/* out0366_em-eta6-phi18*/	7,20,2,4,21,1,6,23,0,1,23,1,3,23,2,16,168,0,15,168,1,3,
/* out0367_em-eta7-phi18*/	5,20,0,2,20,1,13,20,2,8,168,1,13,168,2,3,
/* out0368_em-eta8-phi18*/	7,16,1,1,19,0,5,19,2,8,20,0,1,20,1,3,236,0,2,168,2,13,
/* out0369_em-eta9-phi18*/	6,15,2,5,16,1,1,19,0,11,236,0,9,236,1,2,236,2,13,
/* out0370_em-eta10-phi18*/	6,15,1,10,15,2,3,235,1,8,235,2,5,236,1,1,236,2,3,
/* out0371_em-eta11-phi18*/	6,14,2,6,15,1,5,101,0,7,101,1,3,232,2,2,235,2,11,
/* out0372_em-eta12-phi18*/	6,14,0,7,14,2,2,99,2,1,101,1,11,232,1,6,232,2,4,
/* out0373_em-eta13-phi18*/	7,1,2,2,14,0,5,99,1,5,99,2,6,101,1,1,231,2,3,232,1,7,
/* out0374_em-eta14-phi18*/	6,1,1,5,1,2,2,98,2,1,99,1,8,231,0,2,231,2,5,
/* out0375_em-eta15-phi18*/	5,0,2,1,1,1,5,98,0,2,98,2,7,231,0,6,
/* out0376_em-eta16-phi18*/	5,0,1,1,0,2,4,98,0,6,226,1,3,231,0,2,
/* out0377_em-eta17-phi18*/	6,0,0,2,0,1,1,0,2,3,98,0,3,128,1,2,226,1,4,
/* out0378_em-eta18-phi18*/	4,0,0,5,128,1,4,226,0,2,226,1,2,
/* out0379_em-eta19-phi18*/	2,128,0,2,128,1,2,
/* out0380_em-eta0-phi19*/	1,171,3,10,
/* out0381_em-eta1-phi19*/	2,171,2,12,171,3,6,
/* out0382_em-eta2-phi19*/	2,170,3,14,171,2,4,
/* out0383_em-eta3-phi19*/	2,170,2,15,170,3,2,
/* out0384_em-eta4-phi19*/	2,169,3,16,170,2,1,
/* out0385_em-eta5-phi19*/	9,21,0,1,21,2,12,22,0,8,22,1,16,22,2,6,24,0,1,24,1,7,168,5,1,169,2,16,
/* out0386_em-eta6-phi19*/	7,17,2,2,20,2,1,21,0,12,21,1,10,21,2,2,168,4,3,168,5,15,
/* out0387_em-eta7-phi19*/	7,16,2,1,17,1,8,17,2,1,20,0,11,20,2,3,168,3,3,168,4,13,
/* out0388_em-eta8-phi19*/	8,16,0,1,16,1,5,16,2,11,20,0,2,234,0,2,234,2,1,236,0,2,168,3,13,
/* out0389_em-eta9-phi19*/	7,15,2,5,16,0,1,16,1,9,233,2,1,234,2,5,236,0,3,236,1,11,
/* out0390_em-eta10-phi19*/	5,15,0,10,15,2,3,233,1,6,233,2,9,236,1,2,
/* out0391_em-eta11-phi19*/	8,2,1,1,2,2,4,15,0,5,15,1,1,100,0,10,100,2,3,232,2,4,233,1,9,
/* out0392_em-eta12-phi19*/	8,2,1,7,14,0,3,99,2,2,100,1,1,100,2,12,232,0,5,232,1,1,232,2,6,
/* out0393_em-eta13-phi19*/	8,1,2,6,2,1,1,14,0,1,99,0,4,99,2,7,227,2,1,232,0,6,232,1,2,
/* out0394_em-eta14-phi19*/	9,1,0,1,1,1,1,1,2,4,99,0,7,99,1,2,227,1,4,227,2,1,231,0,3,231,2,1,
/* out0395_em-eta15-phi19*/	10,1,0,2,1,1,4,98,0,2,98,2,1,99,1,1,129,1,3,129,2,2,226,2,1,227,1,3,231,0,3,
/* out0396_em-eta16-phi19*/	7,0,2,3,1,0,1,1,1,1,98,0,3,129,1,3,226,1,4,226,2,1,
/* out0397_em-eta17-phi19*/	5,0,2,4,128,1,4,128,2,2,226,0,2,226,1,3,
/* out0398_em-eta18-phi19*/	5,0,0,3,0,2,1,128,0,1,128,1,4,226,0,4,
/* out0399_em-eta19-phi19*/	1,128,0,5,
/* out0400_em-eta0-phi20*/	1,175,0,10,
/* out0401_em-eta1-phi20*/	2,175,0,6,175,1,12,
/* out0402_em-eta2-phi20*/	2,174,0,14,175,1,4,
/* out0403_em-eta3-phi20*/	2,174,0,2,174,1,15,
/* out0404_em-eta4-phi20*/	3,22,2,1,173,0,16,174,1,1,
/* out0405_em-eta5-phi20*/	8,18,0,1,18,1,3,18,2,14,21,0,1,22,0,8,22,2,9,172,0,1,173,1,16,
/* out0406_em-eta6-phi20*/	7,17,0,1,17,2,10,18,0,2,18,1,13,21,0,2,172,0,15,172,1,3,
/* out0407_em-eta7-phi20*/	6,4,2,1,17,0,12,17,1,7,17,2,3,172,1,13,172,2,3,
/* out0408_em-eta8-phi20*/	8,4,1,5,4,2,2,16,0,8,16,2,4,17,1,1,234,0,10,234,1,1,172,2,13,
/* out0409_em-eta9-phi20*/	7,3,1,1,3,2,9,4,1,1,16,0,6,234,0,3,234,1,7,234,2,10,
/* out0410_em-eta10-phi20*/	7,3,1,11,3,2,1,15,0,1,229,1,1,229,2,1,233,0,8,233,2,6,
/* out0411_em-eta11-phi20*/	9,2,0,1,2,2,10,3,1,1,100,0,6,100,1,6,131,1,2,228,2,4,233,0,8,233,1,1,
/* out0412_em-eta12-phi20*/	9,2,0,4,2,1,4,2,2,1,100,1,9,100,2,1,130,2,3,228,1,7,228,2,1,232,0,3,
/* out0413_em-eta13-phi20*/	10,1,0,1,1,2,2,2,0,1,2,1,3,99,0,3,130,1,6,130,2,2,227,2,6,228,1,2,232,0,2,
/* out0414_em-eta14-phi20*/	7,1,0,6,99,0,2,129,2,5,130,1,3,227,0,1,227,1,3,227,2,4,
/* out0415_em-eta15-phi20*/	5,1,0,5,7,2,1,129,1,2,129,2,5,227,1,6,
/* out0416_em-eta16-phi20*/	4,7,1,1,7,2,3,129,1,6,226,2,6,
/* out0417_em-eta17-phi20*/	5,7,1,4,128,2,5,129,1,1,226,0,3,226,2,3,
/* out0418_em-eta18-phi20*/	4,7,1,2,128,0,2,128,2,4,226,0,3,
/* out0419_em-eta19-phi20*/	1,128,0,4,
/* out0420_em-eta0-phi21*/	1,175,3,10,
/* out0421_em-eta1-phi21*/	2,175,2,12,175,3,6,
/* out0422_em-eta2-phi21*/	2,174,3,14,175,2,4,
/* out0423_em-eta3-phi21*/	2,174,2,15,174,3,2,
/* out0424_em-eta4-phi21*/	2,173,3,16,174,2,1,
/* out0425_em-eta5-phi21*/	6,6,1,9,6,2,9,18,0,6,18,2,2,172,5,1,173,2,16,
/* out0426_em-eta6-phi21*/	7,5,0,1,5,1,4,5,2,14,6,1,3,18,0,7,172,4,3,172,5,15,
/* out0427_em-eta7-phi21*/	6,4,2,8,5,0,1,5,1,12,17,0,3,172,3,3,172,4,13,
/* out0428_em-eta8-phi21*/	8,4,0,7,4,1,7,4,2,5,230,0,3,230,1,5,234,0,1,234,1,3,172,3,13,
/* out0429_em-eta9-phi21*/	8,3,0,4,3,2,6,4,0,1,4,1,3,10,1,1,229,2,8,230,1,7,234,1,5,
/* out0430_em-eta10-phi21*/	6,3,0,10,3,1,2,9,2,1,229,0,1,229,1,11,229,2,4,
/* out0431_em-eta11-phi21*/	11,2,0,3,2,2,1,3,0,1,3,1,1,9,1,3,9,2,2,131,0,5,131,1,7,228,0,1,228,2,9,229,1,3,
/* out0432_em-eta12-phi21*/	8,2,0,6,8,2,2,9,1,2,130,2,8,131,1,7,228,0,5,228,1,4,228,2,2,
/* out0433_em-eta13-phi21*/	10,2,0,1,8,1,1,8,2,6,130,0,5,130,1,3,130,2,3,227,0,1,227,2,3,228,0,1,228,1,3,
/* out0434_em-eta14-phi21*/	6,8,1,6,129,2,3,130,0,2,130,1,4,227,0,7,227,2,1,
/* out0435_em-eta15-phi21*/	6,7,2,4,8,1,2,129,0,7,129,2,1,222,2,1,227,0,5,
/* out0436_em-eta16-phi21*/	5,7,2,4,129,0,6,222,1,2,222,2,1,226,2,2,
/* out0437_em-eta17-phi21*/	9,7,1,4,95,1,2,95,2,2,128,2,1,129,0,1,129,1,1,222,1,2,226,0,1,226,2,3,
/* out0438_em-eta18-phi21*/	4,7,1,3,95,1,2,128,2,3,226,0,1,
/* out0439_em-eta19-phi21*/	2,128,0,2,128,2,1,
/* out0440_em-eta0-phi22*/	1,179,0,10,
/* out0441_em-eta1-phi22*/	2,179,0,6,179,1,12,
/* out0442_em-eta2-phi22*/	2,178,0,14,179,1,4,
/* out0443_em-eta3-phi22*/	2,178,0,2,178,1,15,
/* out0444_em-eta4-phi22*/	2,177,0,16,178,1,1,
/* out0445_em-eta5-phi22*/	8,6,0,14,6,1,2,6,2,7,12,2,3,13,0,2,13,1,8,176,0,1,177,1,16,
/* out0446_em-eta6-phi22*/	8,5,0,7,5,2,2,6,0,2,6,1,2,12,1,9,12,2,5,176,0,15,176,1,3,
/* out0447_em-eta7-phi22*/	6,4,0,1,5,0,7,11,1,4,11,2,11,176,1,13,176,2,3,
/* out0448_em-eta8-phi22*/	5,4,0,7,10,2,5,11,1,8,230,0,7,176,2,13,
/* out0449_em-eta9-phi22*/	9,10,0,1,10,1,8,10,2,8,225,1,3,225,2,4,229,0,2,229,2,3,230,0,6,230,1,4,
/* out0450_em-eta10-phi22*/	6,3,0,1,9,2,7,10,1,5,224,2,2,225,1,2,229,0,12,
/* out0451_em-eta11-phi22*/	10,9,0,2,9,1,4,9,2,5,97,2,1,131,0,7,224,1,5,224,2,4,228,0,2,229,0,1,229,1,1,
/* out0452_em-eta12-phi22*/	9,8,2,3,9,1,6,97,1,4,97,2,5,130,0,2,131,0,4,223,2,3,224,1,3,228,0,6,
/* out0453_em-eta13-phi22*/	8,8,0,2,8,2,5,96,2,2,97,1,4,130,0,6,223,1,3,223,2,6,228,0,1,
/* out0454_em-eta14-phi22*/	7,8,0,3,8,1,4,96,1,2,96,2,7,130,0,1,223,1,6,227,0,1,
/* out0455_em-eta15-phi22*/	6,7,2,2,8,1,3,96,1,7,129,0,1,222,2,6,227,0,1,
/* out0456_em-eta16-phi22*/	7,7,0,3,7,2,2,95,2,5,96,1,1,129,0,1,222,1,3,222,2,3,
/* out0457_em-eta17-phi22*/	4,7,0,4,95,1,2,95,2,4,222,1,5,
/* out0458_em-eta18-phi22*/	4,7,0,2,7,1,1,95,1,5,222,1,1,
/* out0459_em-eta19-phi22*/	2,7,1,1,95,1,1,
/* out0460_em-eta0-phi23*/	1,179,3,10,
/* out0461_em-eta1-phi23*/	2,179,2,12,179,3,6,
/* out0462_em-eta2-phi23*/	2,178,3,14,179,2,4,
/* out0463_em-eta3-phi23*/	2,178,2,15,178,3,2,
/* out0464_em-eta4-phi23*/	2,177,3,16,178,2,1,
/* out0465_em-eta5-phi23*/	6,12,0,1,12,2,5,13,0,14,13,1,8,176,5,1,177,2,16,
/* out0466_em-eta6-phi23*/	5,12,0,15,12,1,6,12,2,3,176,4,3,176,5,15,
/* out0467_em-eta7-phi23*/	5,11,0,11,11,2,5,12,1,1,176,3,3,176,4,13,
/* out0468_em-eta8-phi23*/	7,10,0,1,10,2,2,11,0,5,11,1,4,225,0,7,225,2,3,176,3,13,
/* out0469_em-eta9-phi23*/	5,10,0,12,10,2,1,225,0,7,225,1,4,225,2,9,
/* out0470_em-eta10-phi23*/	8,9,0,2,9,2,1,10,0,2,10,1,2,224,0,7,224,2,6,225,0,2,225,1,7,
/* out0471_em-eta11-phi23*/	6,9,0,9,97,0,1,97,2,5,224,0,7,224,1,3,224,2,4,
/* out0472_em-eta12-phi23*/	9,9,0,3,9,1,1,97,0,13,97,1,2,97,2,5,223,0,1,223,2,4,224,0,2,224,1,5,
/* out0473_em-eta13-phi23*/	8,8,0,5,96,0,1,96,2,3,97,0,2,97,1,6,223,0,6,223,1,1,223,2,3,
/* out0474_em-eta14-phi23*/	5,8,0,5,96,0,5,96,2,4,223,0,3,223,1,5,
/* out0475_em-eta15-phi23*/	7,8,0,1,96,0,4,96,1,5,222,0,2,222,2,4,223,0,6,223,1,1,
/* out0476_em-eta16-phi23*/	7,7,0,3,95,0,7,95,2,4,96,0,6,96,1,1,222,0,5,222,2,1,
/* out0477_em-eta17-phi23*/	5,7,0,3,95,0,5,95,2,1,222,0,3,222,1,2,
/* out0478_em-eta18-phi23*/	5,7,0,1,95,0,3,95,1,2,222,0,6,222,1,1,
/* out0479_em-eta19-phi23*/	2,95,0,1,95,1,2
};