parameter integer matrixH [0:7724] = {
/* num inputs = 235(in0-in234) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 16 */
//* total number of input in adders 2414 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	1,110,0,10,
/* out0002_em-eta2-phi0*/	2,110,0,6,110,1,11,
/* out0003_em-eta3-phi0*/	2,109,0,13,110,1,5,
/* out0004_em-eta4-phi0*/	2,109,0,3,109,1,14,
/* out0005_em-eta5-phi0*/	4,93,1,2,94,1,8,94,2,14,109,1,2,
/* out0006_em-eta6-phi0*/	4,63,2,1,93,0,15,93,1,6,93,2,4,
/* out0007_em-eta7-phi0*/	8,62,0,1,62,1,4,63,1,6,63,2,12,92,0,8,92,1,5,93,0,1,93,2,3,
/* out0008_em-eta8-phi0*/	6,62,0,14,62,1,2,62,2,2,91,1,1,92,0,8,92,2,4,
/* out0009_em-eta9-phi0*/	6,61,0,6,61,1,3,62,0,1,62,2,2,91,0,12,91,1,2,
/* out0010_em-eta10-phi0*/	6,61,0,10,61,2,2,90,0,1,90,1,1,91,0,4,91,2,2,
/* out0011_em-eta11-phi0*/	5,60,0,5,60,1,2,104,0,4,104,1,9,90,0,9,
/* out0012_em-eta12-phi0*/	5,60,0,8,104,0,5,104,1,1,104,2,7,90,0,4,
/* out0013_em-eta13-phi0*/	9,59,0,2,59,1,1,60,0,1,60,2,1,103,0,3,103,1,7,104,0,7,104,2,2,89,0,4,
/* out0014_em-eta14-phi0*/	5,59,0,6,103,0,6,103,1,1,103,2,3,89,0,5,
/* out0015_em-eta15-phi0*/	6,59,0,3,102,0,1,102,1,2,103,0,7,103,2,4,89,0,1,
/* out0016_em-eta16-phi0*/	4,58,0,1,102,0,4,102,1,3,88,0,2,
/* out0017_em-eta17-phi0*/	4,58,0,4,102,0,4,102,2,1,88,0,3,
/* out0018_em-eta18-phi0*/	3,102,0,7,102,2,3,88,0,1,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	1,110,3,10,
/* out0022_em-eta2-phi1*/	2,110,2,11,110,3,6,
/* out0023_em-eta3-phi1*/	2,109,3,13,110,2,5,
/* out0024_em-eta4-phi1*/	2,109,2,14,109,3,3,
/* out0025_em-eta5-phi1*/	7,87,0,12,87,1,7,87,2,1,93,1,1,94,1,8,94,2,2,109,2,2,
/* out0026_em-eta6-phi1*/	9,57,1,1,63,1,1,63,2,2,86,0,5,86,1,3,87,0,4,87,2,3,93,1,7,93,2,7,
/* out0027_em-eta7-phi1*/	9,57,0,13,57,1,1,62,1,4,63,1,9,63,2,1,86,0,10,92,1,11,92,2,1,93,2,2,
/* out0028_em-eta8-phi1*/	7,56,0,4,57,0,1,62,1,6,62,2,10,85,0,7,91,1,3,92,2,11,
/* out0029_em-eta9-phi1*/	6,56,0,4,61,1,12,62,2,2,85,0,1,91,1,10,91,2,5,
/* out0030_em-eta10-phi1*/	6,55,0,1,61,1,1,61,2,13,84,0,1,90,1,5,91,2,8,
/* out0031_em-eta11-phi1*/	6,60,1,11,100,2,10,104,1,6,90,0,2,90,1,7,90,2,3,
/* out0032_em-eta12-phi1*/	6,60,0,2,60,2,8,98,0,5,104,2,7,89,1,2,90,2,8,
/* out0033_em-eta13-phi1*/	6,59,1,6,60,2,2,98,0,4,103,1,6,89,0,2,89,1,7,
/* out0034_em-eta14-phi1*/	7,59,0,3,59,1,2,59,2,1,103,1,2,103,2,6,89,0,3,89,2,3,
/* out0035_em-eta15-phi1*/	8,59,0,2,59,2,5,97,0,1,102,1,2,103,2,3,88,1,2,89,0,1,89,2,3,
/* out0036_em-eta16-phi1*/	5,58,0,2,58,1,4,102,1,6,88,0,3,88,1,2,
/* out0037_em-eta17-phi1*/	4,58,0,5,102,1,1,102,2,5,88,0,4,
/* out0038_em-eta18-phi1*/	3,102,2,3,88,0,3,88,2,1,
/* out0039_em-eta19-phi1*/	1,88,2,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	1,112,0,10,
/* out0042_em-eta2-phi2*/	2,112,0,6,112,1,11,
/* out0043_em-eta3-phi2*/	2,111,0,13,112,1,5,
/* out0044_em-eta4-phi2*/	2,111,0,3,111,1,14,
/* out0045_em-eta5-phi2*/	5,81,0,3,81,1,2,87,1,9,87,2,6,111,1,2,
/* out0046_em-eta6-phi2*/	5,57,1,4,81,0,10,86,1,13,86,2,1,87,2,6,
/* out0047_em-eta7-phi2*/	8,50,0,1,57,0,2,57,1,10,57,2,12,80,0,3,85,1,5,86,0,1,86,2,15,
/* out0048_em-eta8-phi2*/	8,50,0,1,56,0,3,56,1,13,56,2,1,57,2,4,85,0,6,85,1,9,85,2,5,
/* out0049_em-eta9-phi2*/	8,55,1,2,56,0,5,56,2,10,84,0,2,84,1,6,85,0,2,85,2,6,91,2,1,
/* out0050_em-eta10-phi2*/	8,55,0,9,55,1,5,61,2,1,100,1,1,100,2,3,84,0,11,84,1,1,84,2,1,
/* out0051_em-eta11-phi2*/	14,54,1,1,55,0,6,55,2,3,60,1,3,60,2,1,98,1,3,100,1,13,100,2,3,83,0,2,83,1,1,84,0,2,84,2,2,90,1,3,90,2,3,
/* out0052_em-eta12-phi2*/	8,54,0,6,60,2,4,98,0,3,98,1,8,98,2,1,83,0,7,89,1,1,90,2,2,
/* out0053_em-eta13-phi2*/	6,54,0,4,59,1,4,98,0,4,98,2,6,83,0,1,89,1,6,
/* out0054_em-eta14-phi2*/	5,59,1,3,59,2,4,97,0,4,97,1,4,89,2,7,
/* out0055_em-eta15-phi2*/	6,53,0,1,59,2,5,97,0,7,82,0,1,88,1,3,89,2,3,
/* out0056_em-eta16-phi2*/	4,58,1,7,97,0,3,102,1,2,88,1,5,
/* out0057_em-eta17-phi2*/	6,58,0,3,58,1,1,96,1,2,102,2,3,88,1,1,88,2,3,
/* out0058_em-eta18-phi2*/	4,96,0,1,96,1,2,102,2,1,88,2,3,
/* out0059_em-eta19-phi2*/	1,88,2,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	1,112,3,10,
/* out0062_em-eta2-phi3*/	2,112,2,11,112,3,6,
/* out0063_em-eta3-phi3*/	2,111,3,13,112,2,5,
/* out0064_em-eta4-phi3*/	2,111,2,14,111,3,3,
/* out0065_em-eta5-phi3*/	5,76,0,5,76,1,8,76,2,16,81,1,13,111,2,2,
/* out0066_em-eta6-phi3*/	6,52,1,2,75,0,3,80,1,6,81,0,3,81,1,1,81,2,16,
/* out0067_em-eta7-phi3*/	8,50,0,7,50,1,13,50,2,2,52,0,1,52,1,1,80,0,12,80,1,6,80,2,6,
/* out0068_em-eta8-phi3*/	12,49,0,1,49,1,3,50,0,7,50,2,7,56,1,3,56,2,1,79,0,6,79,1,4,80,0,1,80,2,2,85,1,2,85,2,4,
/* out0069_em-eta9-phi3*/	7,49,0,12,49,1,1,55,1,2,56,2,4,79,0,8,84,1,7,85,2,1,
/* out0070_em-eta10-phi3*/	9,49,0,1,55,1,7,55,2,6,100,1,1,101,0,4,101,2,1,78,0,1,84,1,2,84,2,10,
/* out0071_em-eta11-phi3*/	10,48,0,1,54,1,4,55,2,7,100,1,1,101,0,4,101,1,1,101,2,12,78,0,1,83,1,8,84,2,3,
/* out0072_em-eta12-phi3*/	11,54,0,3,54,1,7,54,2,1,98,1,5,98,2,3,99,1,1,101,1,1,101,2,3,83,0,4,83,1,2,83,2,3,
/* out0073_em-eta13-phi3*/	8,54,0,3,54,2,5,97,1,1,98,2,6,99,1,4,82,1,2,83,0,2,83,2,4,
/* out0074_em-eta14-phi3*/	7,53,0,3,53,1,3,54,2,1,59,2,1,97,1,8,82,0,5,82,1,1,
/* out0075_em-eta15-phi3*/	5,53,0,6,97,0,1,97,1,1,97,2,6,82,0,5,
/* out0076_em-eta16-phi3*/	6,53,0,3,58,1,3,96,1,2,97,2,4,82,0,1,88,1,3,
/* out0077_em-eta17-phi3*/	4,58,0,1,58,1,1,96,1,5,88,2,4,
/* out0078_em-eta18-phi3*/	3,96,0,4,96,1,1,88,2,3,
/* out0079_em-eta19-phi3*/	0,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	1,114,0,10,
/* out0082_em-eta2-phi4*/	2,114,0,6,114,1,11,
/* out0083_em-eta3-phi4*/	2,113,0,13,114,1,5,
/* out0084_em-eta4-phi4*/	2,113,0,3,113,1,14,
/* out0085_em-eta5-phi4*/	6,75,1,8,76,0,11,76,1,8,77,0,5,77,1,6,113,1,2,
/* out0086_em-eta6-phi4*/	5,52,1,10,75,0,13,75,1,7,75,2,9,80,1,1,
/* out0087_em-eta7-phi4*/	12,50,1,3,50,2,3,51,1,3,51,2,4,52,0,15,52,1,2,52,2,11,74,0,9,74,1,4,75,2,1,80,1,3,80,2,7,
/* out0088_em-eta8-phi4*/	7,49,1,8,50,2,4,51,1,10,74,0,4,79,1,12,79,2,3,80,2,1,
/* out0089_em-eta9-phi4*/	6,49,0,2,49,1,4,49,2,12,78,1,3,79,0,2,79,2,11,
/* out0090_em-eta10-phi4*/	6,48,0,3,48,1,8,49,2,3,101,0,2,78,0,8,78,1,5,
/* out0091_em-eta11-phi4*/	8,48,0,11,48,2,1,54,1,1,101,0,6,101,1,11,78,0,6,78,2,1,83,1,4,
/* out0092_em-eta12-phi4*/	11,44,1,1,48,0,1,48,2,1,54,1,3,54,2,4,99,1,1,99,2,8,101,1,3,63,1,2,83,1,1,83,2,7,
/* out0093_em-eta13-phi4*/	9,44,1,2,53,1,1,54,2,5,99,0,1,99,1,7,99,2,1,63,1,1,82,1,4,83,2,2,
/* out0094_em-eta14-phi4*/	9,53,1,7,92,1,1,97,1,2,97,2,1,99,0,2,99,1,3,82,0,1,82,1,5,82,2,1,
/* out0095_em-eta15-phi4*/	7,53,0,2,53,1,1,53,2,3,92,1,3,97,2,4,82,0,2,82,2,3,
/* out0096_em-eta16-phi4*/	9,53,0,1,53,2,3,92,1,1,96,1,2,96,2,2,97,2,1,49,1,1,82,0,1,82,2,2,
/* out0097_em-eta17-phi4*/	3,96,1,2,96,2,3,49,1,3,
/* out0098_em-eta18-phi4*/	4,96,0,6,96,2,1,49,0,2,49,1,2,
/* out0099_em-eta19-phi4*/	1,96,0,2,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	1,114,3,10,
/* out0102_em-eta2-phi5*/	2,114,2,11,114,3,6,
/* out0103_em-eta3-phi5*/	2,113,3,13,114,2,5,
/* out0104_em-eta4-phi5*/	2,113,2,14,113,3,3,
/* out0105_em-eta5-phi5*/	5,70,1,2,77,0,11,77,1,10,77,2,16,113,2,2,
/* out0106_em-eta6-phi5*/	9,52,1,1,52,2,1,70,0,3,70,2,3,70,0,14,70,1,5,74,1,1,75,1,1,75,2,6,
/* out0107_em-eta7-phi5*/	10,51,0,2,51,2,12,52,2,4,70,0,2,70,1,8,70,2,13,70,0,2,74,0,1,74,1,11,74,2,10,
/* out0108_em-eta8-phi5*/	8,51,0,14,51,1,3,68,2,4,68,1,3,68,2,8,74,0,2,74,2,6,79,2,1,
/* out0109_em-eta9-phi5*/	6,49,2,1,68,1,12,68,2,4,68,1,13,78,1,2,79,2,1,
/* out0110_em-eta10-phi5*/	5,48,1,8,48,2,2,68,1,4,78,1,6,78,2,8,
/* out0111_em-eta11-phi5*/	7,44,2,1,48,2,11,94,0,9,94,1,1,94,2,10,63,2,4,78,2,7,
/* out0112_em-eta12-phi5*/	8,44,1,2,44,2,7,48,2,1,94,2,6,99,0,1,99,2,6,63,1,6,63,2,3,
/* out0113_em-eta13-phi5*/	5,44,1,9,99,0,9,99,2,1,63,1,7,82,1,1,
/* out0114_em-eta14-phi5*/	7,44,1,2,53,1,4,53,2,1,92,2,5,99,0,3,82,1,3,82,2,4,
/* out0115_em-eta15-phi5*/	4,53,2,6,92,1,5,92,2,2,82,2,5,
/* out0116_em-eta16-phi5*/	5,53,2,3,92,1,6,96,2,1,49,1,3,82,2,1,
/* out0117_em-eta17-phi5*/	2,96,2,5,49,1,4,
/* out0118_em-eta18-phi5*/	4,96,0,1,96,2,4,49,0,4,49,1,1,
/* out0119_em-eta19-phi5*/	1,96,0,2,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	1,116,0,10,
/* out0122_em-eta2-phi6*/	2,116,0,6,116,1,11,
/* out0123_em-eta3-phi6*/	2,115,0,13,116,1,5,
/* out0124_em-eta4-phi6*/	2,115,0,3,115,1,14,
/* out0125_em-eta5-phi6*/	5,70,1,3,72,0,11,72,1,14,72,2,16,115,1,2,
/* out0126_em-eta6-phi6*/	7,70,0,4,71,1,2,69,2,1,70,1,6,70,2,14,71,1,6,71,2,1,
/* out0127_em-eta7-phi6*/	10,69,1,2,69,2,12,70,0,7,70,1,8,71,0,2,71,1,3,69,0,1,69,1,10,69,2,11,70,2,2,
/* out0128_em-eta8-phi6*/	8,68,2,4,69,0,3,69,1,14,65,1,1,68,0,3,68,2,8,69,0,2,69,1,6,
/* out0129_em-eta9-phi6*/	6,46,1,1,68,0,12,68,2,4,64,2,2,65,1,1,68,0,13,
/* out0130_em-eta10-phi6*/	5,45,1,2,45,2,8,68,0,4,64,1,8,64,2,6,
/* out0131_em-eta11-phi6*/	6,44,2,1,45,1,11,94,0,7,94,1,10,63,2,5,64,1,7,
/* out0132_em-eta12-phi6*/	8,44,0,2,44,2,7,45,1,1,93,1,1,93,2,6,94,1,5,63,0,6,63,2,4,
/* out0133_em-eta13-phi6*/	5,44,0,8,93,1,9,93,2,1,50,2,1,63,0,7,
/* out0134_em-eta14-phi6*/	7,39,1,1,39,2,4,44,0,2,92,2,6,93,1,3,50,1,4,50,2,3,
/* out0135_em-eta15-phi6*/	4,39,1,6,92,0,5,92,2,2,50,1,5,
/* out0136_em-eta16-phi6*/	5,39,1,3,92,0,5,49,1,1,49,2,4,50,1,1,
/* out0137_em-eta17-phi6*/	4,105,1,4,49,0,1,49,1,1,49,2,3,
/* out0138_em-eta18-phi6*/	2,105,1,4,49,0,6,
/* out0139_em-eta19-phi6*/	1,105,0,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	1,116,3,10,
/* out0142_em-eta2-phi7*/	2,116,2,11,116,3,6,
/* out0143_em-eta3-phi7*/	2,115,3,13,116,2,5,
/* out0144_em-eta4-phi7*/	2,115,2,14,115,3,3,
/* out0145_em-eta5-phi7*/	7,71,2,8,72,0,5,72,1,2,73,0,16,73,1,12,73,2,2,115,2,2,
/* out0146_em-eta6-phi7*/	6,71,1,8,71,2,3,66,2,1,71,0,13,71,1,9,71,2,7,
/* out0147_em-eta7-phi7*/	12,47,1,3,47,2,3,69,0,3,69,2,4,71,0,14,71,1,3,71,2,10,66,1,7,66,2,3,69,0,9,69,2,4,71,1,1,
/* out0148_em-eta8-phi7*/	7,46,2,8,47,1,4,69,0,10,65,1,3,65,2,12,66,1,1,69,0,4,
/* out0149_em-eta9-phi7*/	6,46,0,2,46,1,12,46,2,4,64,2,3,65,0,2,65,1,11,
/* out0150_em-eta10-phi7*/	6,45,0,3,45,2,8,46,1,3,95,0,2,64,0,8,64,2,5,
/* out0151_em-eta11-phi7*/	9,40,2,1,45,0,11,45,1,1,95,0,8,95,1,1,95,2,11,51,2,4,64,0,6,64,1,1,
/* out0152_em-eta12-phi7*/	11,40,1,4,40,2,3,44,0,2,45,0,1,45,1,1,93,0,1,93,2,8,95,2,4,51,1,7,51,2,1,63,0,2,
/* out0153_em-eta13-phi7*/	9,39,2,1,40,1,5,44,0,2,93,0,7,93,1,1,93,2,1,50,2,4,51,1,2,63,0,1,
/* out0154_em-eta14-phi7*/	10,39,2,7,92,0,1,92,2,1,93,0,3,93,1,2,106,1,1,106,2,2,50,0,1,50,1,1,50,2,5,
/* out0155_em-eta15-phi7*/	7,39,0,2,39,1,3,39,2,1,92,0,3,106,1,4,50,0,2,50,1,3,
/* out0156_em-eta16-phi7*/	9,39,0,1,39,1,3,92,0,2,105,1,2,105,2,1,106,1,1,49,2,2,50,0,1,50,1,2,
/* out0157_em-eta17-phi7*/	3,105,1,4,105,2,1,49,2,5,
/* out0158_em-eta18-phi7*/	4,105,0,5,105,1,2,49,0,3,49,2,2,
/* out0159_em-eta19-phi7*/	1,105,0,2,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	1,118,0,10,
/* out0162_em-eta2-phi8*/	2,118,0,6,118,1,11,
/* out0163_em-eta3-phi8*/	2,117,0,13,118,1,5,
/* out0164_em-eta4-phi8*/	2,117,0,3,117,1,14,
/* out0165_em-eta5-phi8*/	4,67,2,13,73,1,4,73,2,14,117,1,2,
/* out0166_em-eta6-phi8*/	6,71,2,2,66,2,6,67,0,3,67,1,16,67,2,1,71,0,3,
/* out0167_em-eta7-phi8*/	7,47,0,7,47,1,2,47,2,13,71,2,1,66,0,12,66,1,6,66,2,6,
/* out0168_em-eta8-phi8*/	12,42,1,1,42,2,3,46,0,1,46,2,3,47,0,7,47,1,7,53,1,4,53,2,2,65,0,6,65,2,4,66,0,1,66,1,2,
/* out0169_em-eta9-phi8*/	7,41,2,2,42,1,4,46,0,12,46,2,1,52,2,7,53,1,2,65,0,8,
/* out0170_em-eta10-phi8*/	9,41,1,6,41,2,7,46,0,1,95,0,4,95,1,1,108,1,1,52,1,11,52,2,2,64,0,1,
/* out0171_em-eta11-phi8*/	9,40,2,4,41,1,7,45,0,1,95,0,2,95,1,12,108,1,1,51,2,8,52,1,2,64,0,1,
/* out0172_em-eta12-phi8*/	11,40,0,3,40,1,1,40,2,7,93,0,1,95,1,2,95,2,1,107,1,3,107,2,5,51,0,4,51,1,3,51,2,2,
/* out0173_em-eta13-phi8*/	8,40,0,3,40,1,5,93,0,4,106,2,1,107,1,6,50,2,2,51,0,2,51,1,4,
/* out0174_em-eta14-phi8*/	7,34,1,1,39,0,3,39,2,3,40,1,1,106,2,8,50,0,5,50,2,1,
/* out0175_em-eta15-phi8*/	5,39,0,6,106,0,1,106,1,6,106,2,1,50,0,5,
/* out0176_em-eta16-phi8*/	6,33,1,3,39,0,3,105,2,2,106,1,4,50,0,1,56,2,3,
/* out0177_em-eta17-phi8*/	3,33,1,2,105,2,6,56,1,4,
/* out0178_em-eta18-phi8*/	3,105,0,6,105,2,1,56,1,3,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	1,118,3,10,
/* out0182_em-eta2-phi9*/	2,118,2,11,118,3,6,
/* out0183_em-eta3-phi9*/	2,117,3,13,118,2,5,
/* out0184_em-eta4-phi9*/	2,117,2,14,117,3,3,
/* out0185_em-eta5-phi9*/	5,55,1,6,55,2,9,67,0,3,67,2,2,117,2,2,
/* out0186_em-eta6-phi9*/	5,43,2,4,54,1,1,54,2,13,55,1,6,67,0,10,
/* out0187_em-eta7-phi9*/	8,43,0,2,43,1,12,43,2,10,47,0,1,53,2,5,54,0,2,54,1,15,66,0,3,
/* out0188_em-eta8-phi9*/	8,42,0,3,42,1,1,42,2,13,43,1,4,47,0,1,53,0,6,53,1,5,53,2,9,
/* out0189_em-eta9-phi9*/	8,41,2,2,42,0,5,42,1,10,52,0,2,52,2,6,53,0,2,53,1,5,59,1,1,
/* out0190_em-eta10-phi9*/	8,36,1,1,41,0,9,41,2,5,108,0,3,108,1,1,52,0,11,52,1,1,52,2,1,
/* out0191_em-eta11-phi9*/	14,35,1,1,35,2,3,40,2,1,41,0,6,41,1,3,107,2,3,108,0,3,108,1,13,51,0,2,51,2,1,52,0,2,52,1,2,58,1,3,58,2,3,
/* out0192_em-eta12-phi9*/	8,35,1,4,40,0,6,107,0,3,107,1,1,107,2,8,51,0,7,57,2,1,58,1,2,
/* out0193_em-eta13-phi9*/	6,34,2,4,40,0,4,107,0,4,107,1,6,51,0,1,57,2,6,
/* out0194_em-eta14-phi9*/	5,34,1,4,34,2,3,106,0,4,106,2,4,57,1,7,
/* out0195_em-eta15-phi9*/	6,34,1,5,39,0,1,106,0,7,50,0,1,56,2,3,57,1,3,
/* out0196_em-eta16-phi9*/	5,33,1,4,33,2,3,89,2,2,106,0,3,56,2,5,
/* out0197_em-eta17-phi9*/	5,33,1,4,89,1,3,105,2,3,56,1,3,56,2,1,
/* out0198_em-eta18-phi9*/	4,89,1,1,105,0,2,105,2,2,56,1,3,
/* out0199_em-eta19-phi9*/	1,56,1,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	1,120,0,10,
/* out0202_em-eta2-phi10*/	2,120,0,6,120,1,11,
/* out0203_em-eta3-phi10*/	2,119,0,13,120,1,5,
/* out0204_em-eta4-phi10*/	2,119,0,3,119,1,14,
/* out0205_em-eta5-phi10*/	7,55,0,12,55,1,1,55,2,7,61,2,1,62,0,2,62,1,8,119,1,2,
/* out0206_em-eta6-phi10*/	9,38,0,2,38,1,1,43,2,1,54,0,5,54,2,3,55,0,4,55,1,3,61,1,7,61,2,7,
/* out0207_em-eta7-phi10*/	9,37,2,4,38,0,1,38,1,9,43,0,13,43,2,1,54,0,9,60,1,1,60,2,11,61,1,2,
/* out0208_em-eta8-phi10*/	7,37,1,10,37,2,6,42,0,4,43,0,1,53,0,7,59,2,3,60,1,11,
/* out0209_em-eta9-phi10*/	6,36,2,12,37,1,2,42,0,4,53,0,1,59,1,5,59,2,10,
/* out0210_em-eta10-phi10*/	6,36,1,13,36,2,1,41,0,1,52,0,1,58,2,5,59,1,8,
/* out0211_em-eta11-phi10*/	6,35,2,11,91,2,6,108,0,10,58,0,2,58,1,3,58,2,7,
/* out0212_em-eta12-phi10*/	6,35,0,2,35,1,8,91,1,7,107,0,5,57,2,2,58,1,8,
/* out0213_em-eta13-phi10*/	6,34,2,6,35,1,2,90,2,6,107,0,4,57,0,2,57,2,7,
/* out0214_em-eta14-phi10*/	7,34,0,3,34,1,1,34,2,2,90,1,6,90,2,2,57,0,3,57,1,3,
/* out0215_em-eta15-phi10*/	8,34,0,2,34,1,5,89,2,2,90,1,3,106,0,1,56,2,2,57,0,1,57,1,3,
/* out0216_em-eta16-phi10*/	4,33,2,6,89,2,6,56,0,3,56,2,2,
/* out0217_em-eta17-phi10*/	5,33,1,2,33,2,2,89,1,5,89,2,1,56,0,4,
/* out0218_em-eta18-phi10*/	3,89,1,3,56,0,3,56,1,1,
/* out0219_em-eta19-phi10*/	1,56,1,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	1,120,3,10,
/* out0222_em-eta2-phi11*/	2,120,2,11,120,3,6,
/* out0223_em-eta3-phi11*/	2,119,3,13,120,2,5,
/* out0224_em-eta4-phi11*/	2,119,2,14,119,3,3,
/* out0225_em-eta5-phi11*/	5,48,0,5,61,2,2,62,0,14,62,1,8,119,2,2,
/* out0226_em-eta6-phi11*/	6,38,0,1,47,0,1,48,0,3,61,0,15,61,1,4,61,2,6,
/* out0227_em-eta7-phi11*/	10,32,0,6,37,0,1,37,2,4,38,0,12,38,1,6,47,0,6,60,0,8,60,2,5,61,0,1,61,1,3,
/* out0228_em-eta8-phi11*/	9,31,0,2,32,0,1,37,0,14,37,1,2,37,2,2,46,0,5,59,2,1,60,0,8,60,1,4,
/* out0229_em-eta9-phi11*/	8,31,0,6,36,0,6,36,2,3,37,0,1,37,1,2,46,0,2,59,0,12,59,2,2,
/* out0230_em-eta10-phi11*/	8,30,0,3,36,0,10,36,1,2,45,0,6,58,0,1,58,2,1,59,0,4,59,1,2,
/* out0231_em-eta11-phi11*/	7,30,0,5,35,0,5,35,2,2,91,0,4,91,2,9,45,0,2,58,0,9,
/* out0232_em-eta12-phi11*/	7,29,0,2,35,0,8,91,0,5,91,1,7,91,2,1,44,0,4,58,0,4,
/* out0233_em-eta13-phi11*/	10,29,0,5,34,0,2,34,2,1,35,0,1,35,1,1,90,0,2,90,2,7,91,1,2,44,0,3,57,0,4,
/* out0234_em-eta14-phi11*/	7,29,0,1,34,0,6,90,0,5,90,1,3,90,2,1,43,0,1,57,0,5,
/* out0235_em-eta15-phi11*/	7,28,0,3,34,0,3,89,2,2,90,0,1,90,1,4,43,0,4,57,0,1,
/* out0236_em-eta16-phi11*/	6,28,0,4,33,2,2,89,0,3,89,2,3,43,0,3,56,0,2,
/* out0237_em-eta17-phi11*/	6,28,0,1,33,1,1,33,2,3,89,0,4,89,1,1,56,0,3,
/* out0238_em-eta18-phi11*/	4,89,0,1,89,1,3,42,0,3,56,0,1,
/* out0239_em-eta19-phi11*/	2,42,0,1,42,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	1,122,0,10,
/* out0242_em-eta2-phi12*/	2,122,0,6,122,1,11,
/* out0243_em-eta3-phi12*/	2,121,0,13,122,1,5,
/* out0244_em-eta4-phi12*/	2,121,0,3,121,1,14,
/* out0245_em-eta5-phi12*/	5,41,0,2,48,0,5,48,1,15,48,2,2,121,1,2,
/* out0246_em-eta6-phi12*/	6,32,1,1,40,0,1,47,0,2,47,1,10,48,0,3,48,2,13,
/* out0247_em-eta7-phi12*/	6,32,0,7,32,1,13,32,2,5,47,0,7,47,1,4,47,2,13,
/* out0248_em-eta8-phi12*/	7,31,0,2,31,1,10,32,0,2,32,2,8,46,0,6,46,1,12,46,2,2,
/* out0249_em-eta9-phi12*/	6,31,0,6,31,1,2,31,2,9,45,1,4,46,0,3,46,2,9,
/* out0250_em-eta10-phi12*/	6,30,0,3,30,1,9,31,2,2,45,0,6,45,1,6,45,2,2,
/* out0251_em-eta11-phi12*/	9,30,0,5,30,1,1,30,2,7,88,0,11,88,2,1,91,0,3,44,1,3,45,0,2,45,2,7,
/* out0252_em-eta12-phi12*/	9,29,0,2,29,1,6,30,2,2,87,0,6,87,1,2,88,2,1,91,0,4,44,0,5,44,1,5,
/* out0253_em-eta13-phi12*/	7,29,0,5,29,1,1,29,2,3,87,0,8,90,0,2,44,0,4,44,2,4,
/* out0254_em-eta14-phi12*/	11,28,1,2,29,0,1,29,2,4,86,0,2,86,1,1,87,0,1,87,2,1,90,0,5,43,0,1,43,1,4,44,2,2,
/* out0255_em-eta15-phi12*/	6,28,0,3,28,1,3,86,0,6,90,0,1,43,0,4,43,1,1,
/* out0256_em-eta16-phi12*/	6,28,0,4,28,2,1,86,0,3,89,0,3,43,0,3,43,2,2,
/* out0257_em-eta17-phi12*/	6,28,0,1,28,2,3,85,0,2,89,0,4,42,0,3,43,2,2,
/* out0258_em-eta18-phi12*/	4,85,0,3,85,1,1,89,0,1,42,0,4,
/* out0259_em-eta19-phi12*/	1,42,1,2,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	1,122,3,10,
/* out0262_em-eta2-phi13*/	2,122,2,11,122,3,6,
/* out0263_em-eta3-phi13*/	2,121,3,13,122,2,5,
/* out0264_em-eta4-phi13*/	2,121,2,14,121,3,3,
/* out0265_em-eta5-phi13*/	6,40,1,5,41,0,14,41,2,14,48,1,1,48,2,1,121,2,2,
/* out0266_em-eta6-phi13*/	5,27,0,5,40,0,14,40,1,7,40,2,7,47,1,1,
/* out0267_em-eta7-phi13*/	12,26,0,3,26,1,6,27,0,10,27,2,9,32,1,2,32,2,2,39,0,9,39,1,7,40,0,1,40,2,2,47,1,1,47,2,3,
/* out0268_em-eta8-phi13*/	11,26,0,13,26,1,2,26,2,4,31,1,2,32,2,1,38,0,1,38,1,2,39,0,7,39,2,5,46,1,4,46,2,2,
/* out0269_em-eta9-phi13*/	9,25,0,7,25,1,3,26,2,1,31,1,2,31,2,5,38,0,11,38,1,1,45,1,1,46,2,3,
/* out0270_em-eta10-phi13*/	8,25,0,8,25,2,1,30,1,6,37,0,2,38,0,3,38,2,1,45,1,5,45,2,3,
/* out0271_em-eta11-phi13*/	8,24,0,5,30,2,7,84,0,1,88,0,5,88,2,13,37,0,6,44,1,1,45,2,4,
/* out0272_em-eta12-phi13*/	6,24,0,4,29,1,6,87,1,11,37,0,1,44,1,7,44,2,2,
/* out0273_em-eta13-phi13*/	6,29,1,3,29,2,6,87,0,1,87,2,8,36,0,1,44,2,7,
/* out0274_em-eta14-phi13*/	8,23,0,1,28,1,2,29,2,3,86,1,6,87,2,2,36,0,1,43,1,5,44,2,1,
/* out0275_em-eta15-phi13*/	6,28,1,6,86,0,3,86,1,2,86,2,1,43,1,4,43,2,2,
/* out0276_em-eta16-phi13*/	5,28,1,1,28,2,5,86,0,2,86,2,5,43,2,5,
/* out0277_em-eta17-phi13*/	4,28,2,3,85,0,6,42,0,3,43,2,1,
/* out0278_em-eta18-phi13*/	4,85,0,2,85,1,2,42,0,2,42,1,3,
/* out0279_em-eta19-phi13*/	1,42,1,2,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	1,124,0,10,
/* out0282_em-eta2-phi14*/	2,124,0,6,124,1,11,
/* out0283_em-eta3-phi14*/	2,123,0,13,124,1,5,
/* out0284_em-eta4-phi14*/	2,123,0,3,123,1,14,
/* out0285_em-eta5-phi14*/	5,24,0,14,24,1,6,24,2,14,41,2,2,123,1,2,
/* out0286_em-eta6-phi14*/	10,21,0,4,21,2,1,27,0,1,27,2,2,23,0,8,23,1,6,24,1,4,24,2,2,40,1,4,40,2,6,
/* out0287_em-eta7-phi14*/	12,21,0,4,21,1,3,21,2,15,26,1,5,27,2,5,22,0,1,22,1,1,23,0,8,23,2,2,39,1,9,39,2,3,40,2,1,
/* out0288_em-eta8-phi14*/	7,19,0,6,19,1,1,26,1,3,26,2,11,22,0,7,38,1,5,39,2,8,
/* out0289_em-eta9-phi14*/	6,19,0,2,25,1,13,25,2,2,38,0,1,38,1,7,38,2,8,
/* out0290_em-eta10-phi14*/	6,24,1,2,25,0,1,25,2,12,84,1,2,37,1,8,38,2,6,
/* out0291_em-eta11-phi14*/	9,24,0,3,24,1,9,24,2,1,84,0,9,84,1,5,88,2,1,37,0,5,37,1,3,37,2,3,
/* out0292_em-eta12-phi14*/	10,24,0,4,24,2,6,82,1,1,84,0,6,84,2,3,87,1,3,87,2,1,36,1,2,37,0,2,37,2,4,
/* out0293_em-eta13-phi14*/	6,23,0,4,23,1,4,82,0,6,87,2,4,36,0,7,36,1,2,
/* out0294_em-eta14-phi14*/	4,23,0,7,82,0,4,86,1,4,36,0,6,
/* out0295_em-eta15-phi14*/	9,23,0,3,28,1,2,86,1,3,86,2,4,35,0,1,36,0,1,36,2,1,43,1,2,43,2,2,
/* out0296_em-eta16-phi14*/	6,22,1,2,28,2,3,81,0,1,86,2,5,35,0,3,43,2,2,
/* out0297_em-eta17-phi14*/	7,22,0,1,22,1,2,28,2,1,85,0,3,85,1,4,35,0,2,42,1,2,
/* out0298_em-eta18-phi14*/	2,85,1,4,42,1,4,
/* out0299_em-eta19-phi14*/	1,42,1,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	1,124,3,10,
/* out0302_em-eta2-phi15*/	2,124,2,11,124,3,6,
/* out0303_em-eta3-phi15*/	2,123,3,13,124,2,5,
/* out0304_em-eta4-phi15*/	2,123,2,14,123,3,3,
/* out0305_em-eta5-phi15*/	5,24,0,2,24,1,5,28,0,8,28,1,7,123,2,2,
/* out0306_em-eta6-phi15*/	8,21,0,1,23,1,10,23,2,5,24,1,1,26,0,2,26,1,1,28,0,8,28,2,2,
/* out0307_em-eta7-phi15*/	7,19,1,1,20,1,6,21,0,7,21,1,13,22,1,9,23,2,9,26,0,5,
/* out0308_em-eta8-phi15*/	6,19,0,4,19,1,13,19,2,4,22,0,7,22,1,4,22,2,9,
/* out0309_em-eta9-phi15*/	11,17,0,1,17,1,5,19,0,4,19,2,7,25,2,1,21,0,6,21,1,6,22,0,1,22,2,2,38,1,1,38,2,1,
/* out0310_em-eta10-phi15*/	6,17,0,12,17,1,1,84,1,2,21,0,10,21,2,1,37,1,3,
/* out0311_em-eta11-phi15*/	10,16,0,1,17,0,3,17,2,1,24,1,5,24,2,3,84,1,7,84,2,6,20,0,3,37,1,2,37,2,6,
/* out0312_em-eta12-phi15*/	9,16,0,4,23,1,1,24,2,6,82,1,4,83,1,1,84,2,7,20,0,2,36,1,4,37,2,3,
/* out0313_em-eta13-phi15*/	6,23,1,8,82,0,3,82,1,7,82,2,1,36,1,6,36,2,2,
/* out0314_em-eta14-phi15*/	6,23,0,1,23,1,1,23,2,6,82,0,3,82,2,5,36,2,6,
/* out0315_em-eta15-phi15*/	8,22,1,2,23,2,4,81,0,3,81,1,3,82,2,1,86,2,1,35,1,4,36,2,1,
/* out0316_em-eta16-phi15*/	4,22,1,5,81,0,6,35,0,4,35,1,1,
/* out0317_em-eta17-phi15*/	5,22,0,4,22,1,1,81,0,3,85,1,3,35,0,4,
/* out0318_em-eta18-phi15*/	3,85,1,2,35,0,2,42,1,1,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	1,126,0,10,
/* out0322_em-eta2-phi16*/	2,126,0,6,126,1,11,
/* out0323_em-eta3-phi16*/	2,125,0,13,126,1,5,
/* out0324_em-eta4-phi16*/	2,125,0,3,125,1,14,
/* out0325_em-eta5-phi16*/	5,27,1,3,27,2,2,28,1,9,28,2,5,125,1,2,
/* out0326_em-eta6-phi16*/	4,20,2,3,26,1,13,27,1,6,28,2,9,
/* out0327_em-eta7-phi16*/	8,20,0,7,20,1,7,20,2,12,22,1,1,25,1,2,26,0,9,26,1,1,26,2,11,
/* out0328_em-eta8-phi16*/	10,18,1,5,18,2,5,19,1,1,19,2,3,20,0,4,20,1,3,22,1,1,22,2,5,25,0,11,25,1,4,
/* out0329_em-eta9-phi16*/	6,17,1,6,18,1,10,19,2,2,21,1,10,21,2,3,25,0,4,
/* out0330_em-eta10-phi16*/	4,17,1,4,17,2,11,20,1,2,21,2,12,
/* out0331_em-eta11-phi16*/	7,16,0,1,16,1,8,17,2,4,83,1,4,83,2,8,20,0,4,20,1,7,
/* out0332_em-eta12-phi16*/	8,16,0,7,16,1,1,16,2,1,82,1,1,83,0,1,83,1,10,20,0,7,20,2,2,
/* out0333_em-eta13-phi16*/	14,11,1,1,16,0,3,16,2,2,23,1,2,23,2,1,79,0,1,82,1,3,82,2,4,83,0,1,83,1,1,14,1,1,20,2,1,36,1,2,36,2,3,
/* out0334_em-eta14-phi16*/	7,11,1,3,23,2,4,79,0,2,81,1,1,82,2,5,14,1,3,36,2,3,
/* out0335_em-eta15-phi16*/	6,11,1,1,22,1,2,22,2,2,23,2,1,81,1,7,35,1,5,
/* out0336_em-eta16-phi16*/	7,22,1,2,22,2,3,81,0,2,81,1,1,81,2,3,35,1,3,35,2,2,
/* out0337_em-eta17-phi16*/	5,22,0,6,22,2,1,81,0,1,81,2,3,35,2,4,
/* out0338_em-eta18-phi16*/	2,22,0,2,35,2,2,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	1,126,3,10,
/* out0342_em-eta2-phi17*/	2,126,2,11,126,3,6,
/* out0343_em-eta3-phi17*/	2,125,3,13,126,2,5,
/* out0344_em-eta4-phi17*/	2,125,2,14,125,3,3,
/* out0345_em-eta5-phi17*/	4,27,0,3,27,1,1,27,2,14,125,2,2,
/* out0346_em-eta6-phi17*/	6,26,1,1,26,2,1,27,0,13,27,1,6,33,0,1,33,1,6,
/* out0347_em-eta7-phi17*/	8,20,0,4,20,2,1,67,0,10,67,1,7,25,1,3,26,2,4,33,0,15,33,1,1,
/* out0348_em-eta8-phi17*/	7,18,0,4,18,2,11,20,0,1,67,0,6,25,0,1,25,1,7,25,2,11,
/* out0349_em-eta9-phi17*/	6,18,0,12,18,1,1,64,2,4,25,2,5,29,1,2,29,2,7,
/* out0350_em-eta10-phi17*/	4,64,1,10,64,2,4,20,1,1,29,1,12,
/* out0351_em-eta11-phi17*/	8,16,1,6,16,2,1,64,1,6,83,0,2,83,2,8,20,1,6,20,2,5,29,1,1,
/* out0352_em-eta12-phi17*/	6,16,1,1,16,2,9,79,1,1,83,0,11,14,2,1,20,2,8,
/* out0353_em-eta13-phi17*/	7,11,2,5,16,2,3,79,0,3,79,1,7,83,0,1,14,1,2,14,2,6,
/* out0354_em-eta14-phi17*/	4,11,1,5,11,2,2,79,0,8,14,1,7,
/* out0355_em-eta15-phi17*/	7,11,1,6,22,2,1,79,0,2,81,1,4,81,2,1,14,1,3,35,1,2,
/* out0356_em-eta16-phi17*/	4,22,2,5,81,2,6,35,1,1,35,2,4,
/* out0357_em-eta17-phi17*/	4,22,0,1,22,2,4,81,2,3,35,2,4,
/* out0358_em-eta18-phi17*/	1,22,0,2,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	1,128,0,10,
/* out0362_em-eta2-phi18*/	2,128,0,6,128,1,11,
/* out0363_em-eta3-phi18*/	2,127,0,13,128,1,5,
/* out0364_em-eta4-phi18*/	2,127,0,3,127,1,14,
/* out0365_em-eta5-phi18*/	4,34,0,3,34,1,14,34,2,1,127,1,2,
/* out0366_em-eta6-phi18*/	7,67,1,1,31,1,1,31,2,1,33,1,7,33,2,1,34,0,13,34,2,6,
/* out0367_em-eta7-phi18*/	8,66,1,4,66,2,1,67,1,8,67,2,10,30,2,3,31,1,4,33,1,2,33,2,15,
/* out0368_em-eta8-phi18*/	7,65,1,4,65,2,11,66,1,1,67,2,6,30,0,1,30,1,11,30,2,7,
/* out0369_em-eta9-phi18*/	6,64,2,4,65,0,1,65,1,12,29,0,2,29,2,8,30,1,5,
/* out0370_em-eta10-phi18*/	6,64,0,10,64,2,4,15,2,1,29,0,13,29,1,1,29,2,1,
/* out0371_em-eta11-phi18*/	8,12,1,1,12,2,6,64,0,6,80,0,2,80,1,8,15,1,5,15,2,6,29,0,1,
/* out0372_em-eta12-phi18*/	6,12,1,9,12,2,1,79,1,1,80,0,11,14,2,1,15,1,8,
/* out0373_em-eta13-phi18*/	7,11,2,6,12,1,3,79,1,7,79,2,2,80,0,1,14,0,1,14,2,7,
/* out0374_em-eta14-phi18*/	4,11,0,5,11,2,2,79,2,8,14,0,7,
/* out0375_em-eta15-phi18*/	6,11,0,5,76,1,1,76,2,4,79,2,2,7,2,2,14,0,3,
/* out0376_em-eta16-phi18*/	4,5,1,4,76,1,6,7,1,4,7,2,1,
/* out0377_em-eta17-phi18*/	3,5,1,4,76,1,3,7,1,4,
/* out0378_em-eta18-phi18*/	1,5,0,1,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	1,128,3,10,
/* out0382_em-eta2-phi19*/	2,128,2,11,128,3,6,
/* out0383_em-eta3-phi19*/	2,127,3,13,128,2,5,
/* out0384_em-eta4-phi19*/	2,127,2,14,127,3,3,
/* out0385_em-eta5-phi19*/	5,32,1,5,32,2,9,34,1,2,34,2,3,127,2,2,
/* out0386_em-eta6-phi19*/	4,66,2,3,31,2,13,32,1,9,34,2,6,
/* out0387_em-eta7-phi19*/	8,66,0,7,66,1,7,66,2,12,17,2,1,30,2,2,31,0,9,31,1,11,31,2,1,
/* out0388_em-eta8-phi19*/	10,14,1,3,14,2,1,65,0,5,65,2,5,66,0,3,66,1,4,17,1,5,17,2,1,30,0,11,30,2,4,
/* out0389_em-eta9-phi19*/	6,13,2,6,14,1,2,65,0,10,16,1,3,16,2,10,30,0,4,
/* out0390_em-eta10-phi19*/	4,13,1,11,13,2,4,15,2,2,16,1,12,
/* out0391_em-eta11-phi19*/	7,12,0,1,12,2,8,13,1,4,80,1,8,80,2,4,15,0,4,15,2,7,
/* out0392_em-eta12-phi19*/	8,12,0,7,12,1,1,12,2,1,77,2,1,80,0,1,80,2,10,15,0,7,15,1,2,
/* out0393_em-eta13-phi19*/	16,6,1,1,6,2,2,11,0,1,11,2,1,12,0,3,12,1,2,77,1,4,77,2,3,79,2,2,80,0,1,80,2,1,8,1,3,8,2,2,14,0,2,14,2,1,15,1,1,
/* out0394_em-eta14-phi19*/	7,6,1,4,11,0,3,76,2,1,77,1,5,79,2,2,8,1,3,14,0,3,
/* out0395_em-eta15-phi19*/	6,5,1,2,5,2,1,6,1,1,11,0,2,76,2,7,7,2,5,
/* out0396_em-eta16-phi19*/	7,5,1,4,5,2,1,76,0,2,76,1,3,76,2,1,7,1,2,7,2,3,
/* out0397_em-eta17-phi19*/	5,5,0,5,5,1,2,76,0,1,76,1,3,7,1,4,
/* out0398_em-eta18-phi19*/	2,5,0,2,7,1,2,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	1,130,0,10,
/* out0402_em-eta2-phi20*/	2,130,0,6,130,1,11,
/* out0403_em-eta3-phi20*/	2,129,0,13,130,1,5,
/* out0404_em-eta4-phi20*/	2,129,0,3,129,1,14,
/* out0405_em-eta5-phi20*/	5,19,0,3,19,2,6,32,0,8,32,2,7,129,1,2,
/* out0406_em-eta6-phi20*/	8,15,0,1,18,1,5,18,2,10,19,2,2,31,0,2,31,2,1,32,0,8,32,1,2,
/* out0407_em-eta7-phi20*/	8,14,2,1,15,0,9,15,1,1,15,2,15,66,0,6,17,2,9,18,1,9,31,0,5,
/* out0408_em-eta8-phi20*/	6,14,0,4,14,1,4,14,2,13,17,0,7,17,1,9,17,2,4,
/* out0409_em-eta9-phi20*/	11,8,1,1,13,0,1,13,2,5,14,0,4,14,1,7,10,1,1,10,2,1,16,0,6,16,2,6,17,0,1,17,1,2,
/* out0410_em-eta10-phi20*/	6,13,0,12,13,2,1,78,2,2,9,2,3,16,0,10,16,1,1,
/* out0411_em-eta11-phi20*/	10,7,1,3,7,2,5,12,0,1,13,0,3,13,1,1,78,1,6,78,2,7,9,1,6,9,2,2,15,0,3,
/* out0412_em-eta12-phi20*/	9,6,2,1,7,1,6,12,0,4,77,2,4,78,1,7,80,2,1,8,2,4,9,1,3,15,0,2,
/* out0413_em-eta13-phi20*/	6,6,2,8,77,0,3,77,1,1,77,2,7,8,1,2,8,2,6,
/* out0414_em-eta14-phi20*/	6,6,0,1,6,1,6,6,2,1,77,0,3,77,1,5,8,1,6,
/* out0415_em-eta15-phi20*/	8,5,2,2,6,1,4,73,1,1,76,0,3,76,2,3,77,1,1,7,2,4,8,1,1,
/* out0416_em-eta16-phi20*/	4,5,2,6,76,0,6,7,0,4,7,2,1,
/* out0417_em-eta17-phi20*/	5,5,0,6,5,2,1,72,1,3,76,0,3,7,0,4,
/* out0418_em-eta18-phi20*/	3,72,1,2,0,1,2,7,0,2,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	1,130,3,10,
/* out0422_em-eta2-phi21*/	2,130,2,11,130,3,6,
/* out0423_em-eta3-phi21*/	2,129,3,13,130,2,5,
/* out0424_em-eta4-phi21*/	2,129,2,14,129,3,3,
/* out0425_em-eta5-phi21*/	5,13,1,2,19,0,13,19,1,14,19,2,4,129,2,2,
/* out0426_em-eta6-phi21*/	10,10,0,1,10,1,2,15,0,4,15,1,1,12,1,6,12,2,4,18,0,8,18,2,6,19,1,2,19,2,4,
/* out0427_em-eta7-phi21*/	12,9,2,5,10,1,5,15,0,2,15,1,14,15,2,1,11,1,3,11,2,9,12,1,1,17,0,1,17,2,1,18,0,8,18,1,2,
/* out0428_em-eta8-phi21*/	7,9,1,11,9,2,3,14,0,6,14,2,1,10,2,5,11,1,8,17,0,7,
/* out0429_em-eta9-phi21*/	6,8,1,2,8,2,13,14,0,2,10,0,1,10,1,8,10,2,7,
/* out0430_em-eta10-phi21*/	6,7,2,2,8,0,1,8,1,12,78,2,2,9,2,8,10,1,6,
/* out0431_em-eta11-phi21*/	9,7,0,3,7,1,1,7,2,9,75,1,1,78,0,9,78,2,5,9,0,5,9,1,3,9,2,3,
/* out0432_em-eta12-phi21*/	10,7,0,4,7,1,6,74,1,1,74,2,3,77,2,1,78,0,6,78,1,3,8,2,2,9,0,2,9,1,4,
/* out0433_em-eta13-phi21*/	6,6,0,4,6,2,4,74,1,4,77,0,6,8,0,7,8,2,2,
/* out0434_em-eta14-phi21*/	4,6,0,7,73,2,4,77,0,4,8,0,6,
/* out0435_em-eta15-phi21*/	9,0,2,2,6,0,3,73,1,4,73,2,3,1,1,2,1,2,2,7,0,1,8,0,1,8,1,1,
/* out0436_em-eta16-phi21*/	6,0,1,3,5,2,3,73,1,5,76,0,1,1,1,2,7,0,3,
/* out0437_em-eta17-phi21*/	8,0,1,1,5,0,2,5,2,2,72,1,4,72,2,3,0,1,2,0,2,2,7,0,2,
/* out0438_em-eta18-phi21*/	2,72,1,4,0,1,4,
/* out0439_em-eta19-phi21*/	1,0,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	1,132,0,10,
/* out0442_em-eta2-phi22*/	2,132,0,6,132,1,11,
/* out0443_em-eta3-phi22*/	2,131,0,13,132,1,5,
/* out0444_em-eta4-phi22*/	2,131,0,3,131,1,14,
/* out0445_em-eta5-phi22*/	6,6,1,1,6,2,1,12,2,5,13,0,14,13,1,14,131,1,2,
/* out0446_em-eta6-phi22*/	5,10,0,5,5,2,1,12,0,14,12,1,7,12,2,7,
/* out0447_em-eta7-phi22*/	12,4,1,2,4,2,2,9,0,3,9,2,6,10,0,10,10,1,9,5,1,3,5,2,1,11,0,9,11,2,7,12,0,1,12,1,2,
/* out0448_em-eta8-phi22*/	11,3,2,2,4,1,1,9,0,13,9,1,4,9,2,2,4,1,2,4,2,4,10,0,1,10,2,2,11,0,7,11,1,5,
/* out0449_em-eta9-phi22*/	9,3,1,5,3,2,2,8,0,7,8,2,3,9,1,1,3,2,1,4,1,3,10,0,11,10,2,1,
/* out0450_em-eta10-phi22*/	8,2,2,6,8,0,8,8,1,1,3,1,3,3,2,5,9,0,2,10,0,3,10,1,1,
/* out0451_em-eta11-phi22*/	8,2,1,7,7,0,5,75,0,5,75,1,13,78,0,1,2,2,1,3,1,4,9,0,6,
/* out0452_em-eta12-phi22*/	6,1,2,6,7,0,4,74,2,11,2,1,2,2,2,7,9,0,1,
/* out0453_em-eta13-phi22*/	6,1,1,6,1,2,3,74,0,1,74,1,8,2,1,7,8,0,1,
/* out0454_em-eta14-phi22*/	8,0,2,2,1,1,3,6,0,1,73,2,6,74,1,2,1,2,5,2,1,1,8,0,1,
/* out0455_em-eta15-phi22*/	6,0,2,6,73,0,3,73,1,1,73,2,2,1,1,2,1,2,4,
/* out0456_em-eta16-phi22*/	5,0,1,5,0,2,1,73,0,2,73,1,5,1,1,5,
/* out0457_em-eta17-phi22*/	4,0,1,3,72,2,6,0,2,3,1,1,1,
/* out0458_em-eta18-phi22*/	4,72,1,2,72,2,2,0,1,3,0,2,2,
/* out0459_em-eta19-phi22*/	1,0,1,2,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	1,132,3,10,
/* out0462_em-eta2-phi23*/	2,132,2,11,132,3,6,
/* out0463_em-eta3-phi23*/	2,131,3,13,132,2,5,
/* out0464_em-eta4-phi23*/	2,131,2,14,131,3,3,
/* out0465_em-eta5-phi23*/	5,6,0,6,6,1,2,6,2,15,13,0,2,131,2,2,
/* out0466_em-eta6-phi23*/	7,4,0,6,4,2,1,5,0,2,5,2,10,6,0,10,6,1,13,12,0,1,
/* out0467_em-eta7-phi23*/	6,4,0,8,4,1,5,4,2,13,5,0,7,5,1,13,5,2,4,
/* out0468_em-eta8-phi23*/	8,3,0,8,3,2,10,4,0,2,4,1,8,4,0,13,4,1,2,4,2,12,5,0,7,
/* out0469_em-eta9-phi23*/	7,3,0,7,3,1,9,3,2,2,3,0,1,3,2,4,4,0,3,4,1,9,
/* out0470_em-eta10-phi23*/	7,2,0,4,2,2,9,3,0,1,3,1,2,3,0,6,3,1,2,3,2,6,
/* out0471_em-eta11-phi23*/	9,2,0,5,2,1,7,2,2,1,75,0,11,75,1,1,2,0,1,2,2,3,3,0,9,3,1,7,
/* out0472_em-eta12-phi23*/	9,1,0,3,1,2,6,2,0,7,2,1,2,74,0,6,74,2,2,75,1,1,2,0,5,2,2,5,
/* out0473_em-eta13-phi23*/	6,1,0,6,1,1,3,1,2,1,74,0,8,2,0,4,2,1,4,
/* out0474_em-eta14-phi23*/	12,0,0,1,0,2,2,1,0,7,1,1,4,73,0,2,73,2,1,74,0,1,74,1,1,1,0,7,1,2,4,2,0,6,2,1,2,
/* out0475_em-eta15-phi23*/	5,0,0,4,0,2,3,73,0,6,1,0,5,1,2,1,
/* out0476_em-eta16-phi23*/	5,0,0,4,0,1,1,73,0,3,1,0,3,1,1,2,
/* out0477_em-eta17-phi23*/	6,0,0,7,0,1,3,72,2,2,0,2,3,1,0,1,1,1,2,
/* out0478_em-eta18-phi23*/	3,72,1,1,72,2,3,0,2,5,
/* out0479_em-eta19-phi23*/	2,0,1,2,0,2,1
};