parameter integer matrixH [0:6359] = {
/* num inputs = 174(in0-in173) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1933 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	1, 0, 6, 4, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	2, 24, 1, 1, 24, 2, 1, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	2, 3, 5, 4, 3, 11, 7, 
/* out0033_had-eta13-phi1*/	2, 3, 4, 2, 3, 5, 5, 
/* out0034_had-eta14-phi1*/	1, 1, 8, 2, 
/* out0035_had-eta15-phi1*/	3, 1, 5, 1, 1, 8, 1, 1, 11, 12, 
/* out0036_had-eta16-phi1*/	2, 1, 4, 1, 1, 5, 12, 
/* out0037_had-eta17-phi1*/	1, 1, 4, 6, 
/* out0038_had-eta18-phi1*/	1, 0, 3, 6, 
/* out0039_had-eta19-phi1*/	2, 0, 3, 2, 0, 6, 11, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	1, 27, 2, 7, 
/* out0045_had-eta5-phi2*/	3, 26, 2, 1, 27, 1, 12, 27, 2, 4, 
/* out0046_had-eta6-phi2*/	2, 26, 1, 6, 26, 2, 11, 
/* out0047_had-eta7-phi2*/	2, 25, 2, 6, 26, 1, 6, 
/* out0048_had-eta8-phi2*/	2, 25, 1, 9, 25, 2, 5, 
/* out0049_had-eta9-phi2*/	2, 24, 2, 7, 25, 1, 3, 
/* out0050_had-eta10-phi2*/	2, 24, 1, 7, 24, 2, 4, 
/* out0051_had-eta11-phi2*/	3, 3, 8, 13, 3, 9, 2, 24, 1, 4, 
/* out0052_had-eta12-phi2*/	6, 3, 5, 1, 3, 6, 4, 3, 8, 3, 3, 9, 2, 3, 10, 12, 3, 11, 9, 
/* out0053_had-eta13-phi2*/	4, 3, 4, 8, 3, 5, 6, 3, 6, 8, 3, 7, 3, 
/* out0054_had-eta14-phi2*/	4, 1, 8, 11, 1, 9, 2, 3, 4, 6, 3, 7, 1, 
/* out0055_had-eta15-phi2*/	4, 1, 8, 2, 1, 9, 1, 1, 10, 11, 1, 11, 4, 
/* out0056_had-eta16-phi2*/	3, 1, 5, 3, 1, 6, 11, 1, 10, 1, 
/* out0057_had-eta17-phi2*/	2, 1, 4, 8, 1, 7, 3, 
/* out0058_had-eta18-phi2*/	3, 0, 3, 7, 0, 4, 2, 1, 4, 1, 
/* out0059_had-eta19-phi2*/	4, 0, 3, 1, 0, 4, 2, 0, 5, 10, 0, 6, 1, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 118, 0, 5, 
/* out0062_had-eta2-phi3*/	3, 36, 2, 3, 117, 0, 1, 118, 0, 3, 
/* out0063_had-eta3-phi3*/	4, 35, 2, 1, 36, 1, 10, 36, 2, 8, 117, 0, 5, 
/* out0064_had-eta4-phi3*/	6, 27, 0, 4, 27, 2, 4, 35, 1, 7, 35, 2, 8, 116, 0, 2, 117, 0, 2, 
/* out0065_had-eta5-phi3*/	8, 26, 2, 1, 27, 0, 12, 27, 1, 4, 27, 2, 1, 34, 1, 2, 34, 2, 7, 35, 1, 1, 116, 0, 4, 
/* out0066_had-eta6-phi3*/	7, 26, 0, 14, 26, 1, 1, 26, 2, 3, 33, 2, 1, 34, 1, 4, 115, 0, 2, 116, 0, 2, 
/* out0067_had-eta7-phi3*/	7, 25, 0, 3, 25, 2, 4, 26, 0, 2, 26, 1, 3, 33, 1, 3, 33, 2, 3, 115, 0, 3, 
/* out0068_had-eta8-phi3*/	5, 25, 0, 12, 25, 1, 2, 25, 2, 1, 32, 2, 1, 115, 0, 2, 
/* out0069_had-eta9-phi3*/	8, 24, 0, 4, 24, 2, 4, 25, 0, 1, 25, 1, 2, 32, 1, 1, 32, 2, 1, 114, 0, 3, 115, 0, 1, 
/* out0070_had-eta10-phi3*/	3, 24, 0, 9, 24, 1, 1, 114, 0, 5, 
/* out0071_had-eta11-phi3*/	4, 3, 3, 5, 3, 9, 10, 24, 0, 1, 24, 1, 3, 
/* out0072_had-eta12-phi3*/	6, 3, 0, 1, 3, 1, 1, 3, 2, 11, 3, 3, 9, 3, 9, 2, 3, 10, 4, 
/* out0073_had-eta13-phi3*/	4, 3, 1, 10, 3, 2, 5, 3, 6, 4, 3, 7, 6, 
/* out0074_had-eta14-phi3*/	4, 1, 3, 3, 1, 9, 11, 3, 1, 1, 3, 7, 6, 
/* out0075_had-eta15-phi3*/	4, 1, 2, 7, 1, 3, 4, 1, 9, 2, 1, 10, 4, 
/* out0076_had-eta16-phi3*/	3, 1, 1, 2, 1, 2, 9, 1, 6, 4, 
/* out0077_had-eta17-phi3*/	3, 1, 1, 1, 1, 6, 1, 1, 7, 11, 
/* out0078_had-eta18-phi3*/	2, 0, 4, 9, 1, 7, 1, 
/* out0079_had-eta19-phi3*/	4, 0, 1, 14, 0, 2, 1, 0, 4, 2, 0, 5, 6, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 118, 0, 5, 
/* out0082_had-eta2-phi4*/	4, 36, 0, 2, 36, 2, 3, 117, 0, 1, 118, 0, 3, 
/* out0083_had-eta3-phi4*/	8, 35, 0, 1, 35, 2, 2, 36, 0, 14, 36, 1, 6, 36, 2, 2, 46, 1, 3, 46, 2, 9, 117, 0, 5, 
/* out0084_had-eta4-phi4*/	7, 35, 0, 15, 35, 1, 6, 35, 2, 5, 45, 2, 4, 46, 1, 4, 116, 0, 2, 117, 0, 2, 
/* out0085_had-eta5-phi4*/	7, 34, 0, 11, 34, 1, 1, 34, 2, 9, 35, 1, 2, 45, 1, 2, 45, 2, 1, 116, 0, 4, 
/* out0086_had-eta6-phi4*/	6, 33, 0, 2, 33, 2, 7, 34, 0, 4, 34, 1, 9, 115, 0, 2, 116, 0, 2, 
/* out0087_had-eta7-phi4*/	4, 33, 0, 6, 33, 1, 9, 33, 2, 5, 115, 0, 3, 
/* out0088_had-eta8-phi4*/	3, 32, 2, 11, 33, 1, 4, 115, 0, 2, 
/* out0089_had-eta9-phi4*/	5, 32, 0, 1, 32, 1, 10, 32, 2, 2, 114, 0, 3, 115, 0, 1, 
/* out0090_had-eta10-phi4*/	4, 5, 2, 7, 24, 0, 2, 32, 1, 2, 114, 0, 5, 
/* out0091_had-eta11-phi4*/	2, 5, 1, 5, 5, 2, 4, 
/* out0092_had-eta12-phi4*/	4, 3, 0, 11, 3, 3, 2, 4, 8, 3, 5, 1, 4, 
/* out0093_had-eta13-phi4*/	4, 3, 0, 4, 3, 1, 4, 4, 8, 7, 4, 11, 10, 
/* out0094_had-eta14-phi4*/	3, 1, 3, 3, 4, 5, 13, 4, 11, 5, 
/* out0095_had-eta15-phi4*/	3, 1, 0, 8, 1, 3, 6, 4, 4, 3, 
/* out0096_had-eta16-phi4*/	3, 1, 0, 7, 1, 1, 7, 2, 8, 1, 
/* out0097_had-eta17-phi4*/	3, 1, 1, 6, 1, 7, 1, 2, 11, 5, 
/* out0098_had-eta18-phi4*/	3, 0, 2, 6, 0, 4, 1, 2, 5, 3, 
/* out0099_had-eta19-phi4*/	3, 0, 0, 1, 0, 1, 2, 0, 2, 8, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 123, 0, 5, 
/* out0102_had-eta2-phi5*/	2, 122, 0, 1, 123, 0, 3, 
/* out0103_had-eta3-phi5*/	6, 46, 0, 14, 46, 1, 2, 46, 2, 7, 55, 2, 3, 56, 1, 9, 122, 0, 5, 
/* out0104_had-eta4-phi5*/	8, 45, 0, 9, 45, 2, 11, 46, 0, 2, 46, 1, 7, 55, 1, 2, 55, 2, 2, 121, 0, 2, 122, 0, 2, 
/* out0105_had-eta5-phi5*/	6, 34, 0, 1, 44, 0, 1, 44, 2, 8, 45, 0, 4, 45, 1, 14, 121, 0, 4, 
/* out0106_had-eta6-phi5*/	6, 33, 0, 1, 44, 0, 2, 44, 1, 12, 44, 2, 8, 120, 0, 2, 121, 0, 2, 
/* out0107_had-eta7-phi5*/	4, 33, 0, 7, 43, 2, 10, 44, 1, 2, 120, 0, 3, 
/* out0108_had-eta8-phi5*/	5, 32, 0, 7, 32, 2, 1, 43, 1, 7, 43, 2, 1, 120, 0, 2, 
/* out0109_had-eta9-phi5*/	5, 32, 0, 8, 32, 1, 2, 42, 2, 3, 119, 0, 3, 120, 0, 1, 
/* out0110_had-eta10-phi5*/	5, 5, 0, 5, 5, 2, 4, 32, 1, 1, 42, 1, 1, 119, 0, 5, 
/* out0111_had-eta11-phi5*/	3, 5, 0, 5, 5, 1, 3, 5, 2, 1, 
/* out0112_had-eta12-phi5*/	3, 4, 8, 4, 4, 9, 9, 5, 1, 4, 
/* out0113_had-eta13-phi5*/	5, 4, 2, 2, 4, 8, 2, 4, 9, 5, 4, 10, 14, 4, 11, 1, 
/* out0114_had-eta14-phi5*/	6, 4, 2, 1, 4, 4, 1, 4, 5, 3, 4, 6, 13, 4, 7, 1, 4, 10, 2, 
/* out0115_had-eta15-phi5*/	4, 1, 0, 1, 2, 8, 3, 4, 4, 12, 4, 7, 2, 
/* out0116_had-eta16-phi5*/	2, 2, 8, 11, 2, 11, 3, 
/* out0117_had-eta17-phi5*/	4, 2, 5, 1, 2, 6, 1, 2, 10, 3, 2, 11, 8, 
/* out0118_had-eta18-phi5*/	1, 2, 5, 10, 
/* out0119_had-eta19-phi5*/	3, 0, 0, 15, 0, 2, 1, 2, 4, 4, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 123, 0, 5, 
/* out0122_had-eta2-phi6*/	4, 56, 0, 4, 108, 2, 3, 122, 0, 1, 123, 0, 3, 
/* out0123_had-eta3-phi6*/	7, 55, 0, 8, 55, 2, 9, 56, 0, 12, 56, 1, 7, 108, 1, 5, 108, 2, 8, 122, 0, 5, 
/* out0124_had-eta4-phi6*/	8, 45, 0, 2, 54, 0, 1, 54, 2, 7, 55, 0, 7, 55, 1, 14, 55, 2, 2, 121, 0, 2, 122, 0, 2, 
/* out0125_had-eta5-phi6*/	6, 44, 0, 3, 45, 0, 1, 54, 0, 2, 54, 1, 12, 54, 2, 9, 121, 0, 4, 
/* out0126_had-eta6-phi6*/	7, 44, 0, 10, 44, 1, 2, 53, 1, 2, 53, 2, 8, 54, 1, 1, 120, 0, 2, 121, 0, 2, 
/* out0127_had-eta7-phi6*/	4, 43, 0, 10, 43, 2, 5, 53, 1, 2, 120, 0, 3, 
/* out0128_had-eta8-phi6*/	4, 42, 2, 3, 43, 0, 3, 43, 1, 9, 120, 0, 2, 
/* out0129_had-eta9-phi6*/	5, 42, 0, 1, 42, 1, 2, 42, 2, 10, 119, 0, 3, 120, 0, 1, 
/* out0130_had-eta10-phi6*/	4, 5, 0, 1, 6, 8, 2, 42, 1, 9, 119, 0, 5, 
/* out0131_had-eta11-phi6*/	3, 5, 0, 4, 6, 8, 11, 6, 11, 9, 
/* out0132_had-eta12-phi6*/	6, 4, 3, 7, 4, 9, 2, 5, 0, 1, 6, 4, 1, 6, 5, 10, 6, 11, 6, 
/* out0133_had-eta13-phi6*/	4, 4, 0, 6, 4, 1, 1, 4, 2, 8, 4, 3, 9, 
/* out0134_had-eta14-phi6*/	4, 4, 1, 9, 4, 2, 5, 4, 6, 3, 4, 7, 4, 
/* out0135_had-eta15-phi6*/	3, 2, 8, 1, 2, 9, 7, 4, 7, 9, 
/* out0136_had-eta16-phi6*/	2, 2, 9, 7, 2, 10, 7, 
/* out0137_had-eta17-phi6*/	3, 2, 2, 1, 2, 6, 5, 2, 10, 6, 
/* out0138_had-eta18-phi6*/	4, 2, 4, 1, 2, 5, 2, 2, 6, 6, 2, 7, 1, 
/* out0139_had-eta19-phi6*/	1, 2, 4, 9, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 128, 0, 5, 
/* out0142_had-eta2-phi7*/	5, 108, 0, 2, 108, 2, 2, 109, 2, 1, 127, 0, 1, 128, 0, 3, 
/* out0143_had-eta3-phi7*/	9, 55, 0, 1, 107, 0, 3, 107, 2, 6, 108, 0, 14, 108, 1, 11, 108, 2, 3, 109, 1, 1, 109, 2, 5, 127, 0, 5, 
/* out0144_had-eta4-phi7*/	7, 54, 0, 3, 106, 2, 1, 107, 0, 5, 107, 1, 14, 107, 2, 10, 126, 0, 2, 127, 0, 2, 
/* out0145_had-eta5-phi7*/	7, 53, 0, 1, 53, 2, 1, 54, 0, 10, 54, 1, 3, 106, 1, 3, 106, 2, 9, 126, 0, 4, 
/* out0146_had-eta6-phi7*/	6, 53, 0, 12, 53, 1, 4, 53, 2, 7, 106, 1, 1, 125, 0, 2, 126, 0, 2, 
/* out0147_had-eta7-phi7*/	4, 43, 0, 2, 52, 2, 9, 53, 1, 8, 125, 0, 3, 
/* out0148_had-eta8-phi7*/	5, 42, 0, 2, 43, 0, 1, 52, 1, 7, 52, 2, 6, 125, 0, 2, 
/* out0149_had-eta9-phi7*/	4, 42, 0, 11, 52, 1, 1, 124, 0, 3, 125, 0, 1, 
/* out0150_had-eta10-phi7*/	7, 6, 3, 4, 6, 8, 1, 6, 9, 9, 42, 0, 2, 42, 1, 4, 62, 2, 1, 124, 0, 5, 
/* out0151_had-eta11-phi7*/	7, 6, 2, 8, 6, 3, 2, 6, 6, 1, 6, 8, 2, 6, 9, 7, 6, 10, 15, 6, 11, 1, 
/* out0152_had-eta12-phi7*/	5, 6, 4, 6, 6, 5, 6, 6, 6, 14, 6, 7, 3, 6, 10, 1, 
/* out0153_had-eta13-phi7*/	3, 4, 0, 8, 6, 4, 8, 7, 8, 7, 
/* out0154_had-eta14-phi7*/	4, 4, 0, 2, 4, 1, 5, 7, 8, 3, 7, 11, 10, 
/* out0155_had-eta15-phi7*/	5, 2, 3, 6, 2, 9, 2, 4, 1, 1, 7, 5, 6, 7, 11, 2, 
/* out0156_had-eta16-phi7*/	2, 2, 2, 4, 2, 3, 10, 
/* out0157_had-eta17-phi7*/	3, 2, 1, 1, 2, 2, 10, 2, 6, 1, 
/* out0158_had-eta18-phi7*/	4, 2, 1, 1, 2, 2, 1, 2, 6, 3, 2, 7, 6, 
/* out0159_had-eta19-phi7*/	2, 2, 4, 2, 2, 7, 4, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 128, 0, 5, 
/* out0162_had-eta2-phi8*/	4, 109, 0, 2, 109, 2, 3, 127, 0, 1, 128, 0, 3, 
/* out0163_had-eta3-phi8*/	6, 96, 2, 4, 107, 0, 1, 109, 0, 14, 109, 1, 15, 109, 2, 7, 127, 0, 5, 
/* out0164_had-eta4-phi8*/	8, 96, 1, 7, 96, 2, 12, 106, 0, 2, 106, 2, 2, 107, 0, 7, 107, 1, 2, 126, 0, 2, 127, 0, 2, 
/* out0165_had-eta5-phi8*/	4, 106, 0, 14, 106, 1, 9, 106, 2, 4, 126, 0, 4, 
/* out0166_had-eta6-phi8*/	6, 53, 0, 3, 94, 1, 1, 94, 2, 15, 106, 1, 3, 125, 0, 2, 126, 0, 2, 
/* out0167_had-eta7-phi8*/	5, 52, 0, 9, 52, 2, 1, 94, 1, 7, 94, 2, 1, 125, 0, 3, 
/* out0168_had-eta8-phi8*/	4, 52, 0, 7, 52, 1, 7, 62, 2, 1, 125, 0, 2, 
/* out0169_had-eta9-phi8*/	4, 52, 1, 1, 62, 2, 12, 124, 0, 3, 125, 0, 1, 
/* out0170_had-eta10-phi8*/	4, 6, 3, 4, 62, 1, 7, 62, 2, 2, 124, 0, 5, 
/* out0171_had-eta11-phi8*/	4, 6, 0, 16, 6, 1, 5, 6, 2, 6, 6, 3, 6, 
/* out0172_had-eta12-phi8*/	5, 6, 1, 11, 6, 2, 2, 6, 6, 1, 6, 7, 12, 7, 9, 1, 
/* out0173_had-eta13-phi8*/	5, 6, 4, 1, 6, 7, 1, 7, 8, 6, 7, 9, 14, 7, 10, 4, 
/* out0174_had-eta14-phi8*/	3, 7, 6, 5, 7, 10, 11, 7, 11, 4, 
/* out0175_had-eta15-phi8*/	3, 7, 4, 4, 7, 5, 10, 7, 6, 2, 
/* out0176_had-eta16-phi8*/	2, 2, 0, 11, 7, 4, 3, 
/* out0177_had-eta17-phi8*/	2, 2, 0, 5, 2, 1, 7, 
/* out0178_had-eta18-phi8*/	2, 2, 1, 7, 2, 7, 3, 
/* out0179_had-eta19-phi8*/	1, 2, 7, 2, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 133, 0, 5, 
/* out0182_had-eta2-phi9*/	4, 98, 0, 3, 98, 2, 2, 132, 0, 1, 133, 0, 3, 
/* out0183_had-eta3-phi9*/	6, 96, 0, 4, 97, 2, 1, 98, 0, 7, 98, 1, 15, 98, 2, 14, 132, 0, 5, 
/* out0184_had-eta4-phi9*/	8, 95, 0, 2, 95, 2, 2, 96, 0, 12, 96, 1, 8, 97, 1, 2, 97, 2, 7, 131, 0, 2, 132, 0, 2, 
/* out0185_had-eta5-phi9*/	5, 95, 0, 4, 95, 1, 9, 95, 2, 14, 96, 1, 1, 131, 0, 4, 
/* out0186_had-eta6-phi9*/	6, 64, 2, 3, 94, 0, 15, 94, 1, 1, 95, 1, 3, 130, 0, 2, 131, 0, 2, 
/* out0187_had-eta7-phi9*/	5, 63, 0, 1, 63, 2, 9, 94, 0, 1, 94, 1, 7, 130, 0, 3, 
/* out0188_had-eta8-phi9*/	4, 62, 0, 1, 63, 1, 7, 63, 2, 7, 130, 0, 2, 
/* out0189_had-eta9-phi9*/	4, 62, 0, 11, 63, 1, 1, 129, 0, 3, 130, 0, 1, 
/* out0190_had-eta10-phi9*/	4, 8, 9, 4, 62, 0, 2, 62, 1, 8, 129, 0, 5, 
/* out0191_had-eta11-phi9*/	5, 8, 8, 16, 8, 9, 6, 8, 10, 6, 8, 11, 5, 62, 1, 1, 
/* out0192_had-eta12-phi9*/	5, 7, 3, 2, 8, 5, 12, 8, 6, 1, 8, 10, 2, 8, 11, 11, 
/* out0193_had-eta13-phi9*/	6, 7, 0, 4, 7, 2, 4, 7, 3, 14, 7, 9, 1, 8, 4, 1, 8, 5, 1, 
/* out0194_had-eta14-phi9*/	4, 7, 1, 3, 7, 2, 12, 7, 6, 6, 7, 10, 1, 
/* out0195_had-eta15-phi9*/	3, 7, 4, 5, 7, 6, 3, 7, 7, 9, 
/* out0196_had-eta16-phi9*/	2, 7, 4, 4, 9, 8, 11, 
/* out0197_had-eta17-phi9*/	2, 9, 8, 5, 9, 11, 7, 
/* out0198_had-eta18-phi9*/	2, 9, 5, 3, 9, 11, 7, 
/* out0199_had-eta19-phi9*/	1, 9, 5, 2, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 133, 0, 5, 
/* out0202_had-eta2-phi10*/	5, 98, 0, 1, 99, 0, 2, 99, 2, 2, 132, 0, 1, 133, 0, 3, 
/* out0203_had-eta3-phi10*/	9, 66, 2, 1, 97, 0, 6, 97, 2, 3, 98, 0, 5, 98, 1, 1, 99, 0, 3, 99, 1, 11, 99, 2, 14, 132, 0, 5, 
/* out0204_had-eta4-phi10*/	7, 65, 2, 3, 95, 0, 1, 97, 0, 10, 97, 1, 14, 97, 2, 5, 131, 0, 2, 132, 0, 2, 
/* out0205_had-eta5-phi10*/	7, 64, 0, 1, 64, 2, 1, 65, 1, 3, 65, 2, 10, 95, 0, 9, 95, 1, 3, 131, 0, 4, 
/* out0206_had-eta6-phi10*/	6, 64, 0, 7, 64, 1, 4, 64, 2, 12, 95, 1, 1, 130, 0, 2, 131, 0, 2, 
/* out0207_had-eta7-phi10*/	4, 63, 0, 9, 64, 1, 8, 75, 2, 2, 130, 0, 3, 
/* out0208_had-eta8-phi10*/	5, 63, 0, 6, 63, 1, 7, 74, 2, 2, 75, 2, 1, 130, 0, 2, 
/* out0209_had-eta9-phi10*/	5, 62, 0, 1, 63, 1, 1, 74, 2, 11, 129, 0, 3, 130, 0, 1, 
/* out0210_had-eta10-phi10*/	7, 8, 0, 1, 8, 3, 9, 8, 9, 4, 62, 0, 1, 74, 1, 4, 74, 2, 2, 129, 0, 5, 
/* out0211_had-eta11-phi10*/	7, 8, 0, 2, 8, 1, 1, 8, 2, 15, 8, 3, 7, 8, 6, 1, 8, 9, 2, 8, 10, 8, 
/* out0212_had-eta12-phi10*/	5, 8, 2, 1, 8, 4, 6, 8, 5, 3, 8, 6, 14, 8, 7, 6, 
/* out0213_had-eta13-phi10*/	3, 7, 0, 9, 8, 4, 8, 10, 8, 8, 
/* out0214_had-eta14-phi10*/	4, 7, 0, 3, 7, 1, 11, 10, 8, 2, 10, 11, 5, 
/* out0215_had-eta15-phi10*/	5, 7, 1, 2, 7, 7, 7, 9, 3, 2, 9, 9, 6, 10, 11, 1, 
/* out0216_had-eta16-phi10*/	2, 9, 9, 10, 9, 10, 4, 
/* out0217_had-eta17-phi10*/	3, 9, 6, 1, 9, 10, 10, 9, 11, 1, 
/* out0218_had-eta18-phi10*/	4, 9, 5, 6, 9, 6, 3, 9, 10, 1, 9, 11, 1, 
/* out0219_had-eta19-phi10*/	2, 9, 4, 2, 9, 5, 4, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 138, 0, 5, 
/* out0222_had-eta2-phi11*/	4, 67, 1, 4, 99, 0, 3, 137, 0, 1, 138, 0, 3, 
/* out0223_had-eta3-phi11*/	7, 66, 0, 9, 66, 2, 8, 67, 0, 7, 67, 1, 12, 99, 0, 8, 99, 1, 5, 137, 0, 5, 
/* out0224_had-eta4-phi11*/	8, 65, 0, 7, 65, 2, 1, 66, 0, 2, 66, 1, 14, 66, 2, 7, 77, 2, 2, 136, 0, 2, 137, 0, 2, 
/* out0225_had-eta5-phi11*/	6, 65, 0, 9, 65, 1, 12, 65, 2, 2, 76, 2, 3, 77, 2, 1, 136, 0, 4, 
/* out0226_had-eta6-phi11*/	7, 64, 0, 8, 64, 1, 2, 65, 1, 1, 76, 1, 2, 76, 2, 10, 135, 0, 2, 136, 0, 2, 
/* out0227_had-eta7-phi11*/	4, 64, 1, 2, 75, 0, 5, 75, 2, 10, 135, 0, 3, 
/* out0228_had-eta8-phi11*/	4, 74, 0, 3, 75, 1, 9, 75, 2, 3, 135, 0, 2, 
/* out0229_had-eta9-phi11*/	5, 74, 0, 10, 74, 1, 2, 74, 2, 1, 134, 0, 3, 135, 0, 1, 
/* out0230_had-eta10-phi11*/	4, 8, 0, 2, 11, 2, 1, 74, 1, 9, 134, 0, 5, 
/* out0231_had-eta11-phi11*/	3, 8, 0, 11, 8, 1, 9, 11, 2, 4, 
/* out0232_had-eta12-phi11*/	6, 8, 1, 6, 8, 4, 1, 8, 7, 10, 10, 3, 2, 10, 9, 7, 11, 2, 1, 
/* out0233_had-eta13-phi11*/	4, 10, 8, 6, 10, 9, 9, 10, 10, 8, 10, 11, 1, 
/* out0234_had-eta14-phi11*/	4, 10, 5, 4, 10, 6, 3, 10, 10, 5, 10, 11, 9, 
/* out0235_had-eta15-phi11*/	3, 9, 0, 1, 9, 3, 7, 10, 5, 9, 
/* out0236_had-eta16-phi11*/	2, 9, 2, 7, 9, 3, 7, 
/* out0237_had-eta17-phi11*/	3, 9, 2, 6, 9, 6, 5, 9, 10, 1, 
/* out0238_had-eta18-phi11*/	4, 9, 4, 2, 9, 5, 1, 9, 6, 6, 9, 7, 2, 
/* out0239_had-eta19-phi11*/	1, 9, 4, 8, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 138, 0, 5, 
/* out0242_had-eta2-phi12*/	2, 137, 0, 1, 138, 0, 3, 
/* out0243_had-eta3-phi12*/	6, 66, 0, 3, 67, 0, 9, 78, 0, 7, 78, 1, 2, 78, 2, 14, 137, 0, 5, 
/* out0244_had-eta4-phi12*/	8, 66, 0, 2, 66, 1, 2, 77, 0, 11, 77, 2, 9, 78, 1, 7, 78, 2, 2, 136, 0, 2, 137, 0, 2, 
/* out0245_had-eta5-phi12*/	6, 76, 0, 8, 76, 2, 1, 77, 1, 14, 77, 2, 4, 86, 2, 1, 136, 0, 4, 
/* out0246_had-eta6-phi12*/	6, 76, 0, 8, 76, 1, 12, 76, 2, 2, 85, 2, 1, 135, 0, 2, 136, 0, 2, 
/* out0247_had-eta7-phi12*/	4, 75, 0, 10, 76, 1, 2, 85, 2, 7, 135, 0, 3, 
/* out0248_had-eta8-phi12*/	5, 75, 0, 1, 75, 1, 7, 84, 0, 1, 84, 2, 7, 135, 0, 2, 
/* out0249_had-eta9-phi12*/	5, 74, 0, 3, 84, 1, 2, 84, 2, 8, 134, 0, 3, 135, 0, 1, 
/* out0250_had-eta10-phi12*/	5, 11, 0, 4, 11, 2, 5, 74, 1, 1, 84, 1, 1, 134, 0, 5, 
/* out0251_had-eta11-phi12*/	3, 11, 0, 1, 11, 1, 3, 11, 2, 5, 
/* out0252_had-eta12-phi12*/	3, 10, 0, 4, 10, 3, 9, 11, 1, 4, 
/* out0253_had-eta13-phi12*/	5, 10, 0, 2, 10, 1, 1, 10, 2, 14, 10, 3, 5, 10, 10, 2, 
/* out0254_had-eta14-phi12*/	6, 10, 2, 2, 10, 4, 1, 10, 5, 1, 10, 6, 13, 10, 7, 3, 10, 10, 1, 
/* out0255_had-eta15-phi12*/	3, 9, 0, 3, 10, 4, 12, 10, 5, 2, 
/* out0256_had-eta16-phi12*/	2, 9, 0, 11, 9, 1, 3, 
/* out0257_had-eta17-phi12*/	4, 9, 1, 8, 9, 2, 3, 9, 6, 1, 9, 7, 1, 
/* out0258_had-eta18-phi12*/	1, 9, 7, 10, 
/* out0259_had-eta19-phi12*/	2, 9, 4, 4, 12, 4, 14, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 143, 0, 5, 
/* out0262_had-eta2-phi13*/	4, 88, 0, 3, 88, 2, 2, 142, 0, 1, 143, 0, 3, 
/* out0263_had-eta3-phi13*/	8, 78, 0, 9, 78, 1, 3, 87, 0, 2, 87, 2, 1, 88, 0, 2, 88, 1, 6, 88, 2, 14, 142, 0, 5, 
/* out0264_had-eta4-phi13*/	7, 77, 0, 4, 78, 1, 4, 87, 0, 5, 87, 1, 6, 87, 2, 15, 141, 0, 2, 142, 0, 2, 
/* out0265_had-eta5-phi13*/	7, 77, 0, 1, 77, 1, 2, 86, 0, 9, 86, 1, 1, 86, 2, 11, 87, 1, 2, 141, 0, 4, 
/* out0266_had-eta6-phi13*/	6, 85, 0, 7, 85, 2, 2, 86, 1, 9, 86, 2, 4, 140, 0, 2, 141, 0, 2, 
/* out0267_had-eta7-phi13*/	4, 85, 0, 5, 85, 1, 9, 85, 2, 6, 140, 0, 3, 
/* out0268_had-eta8-phi13*/	3, 84, 0, 11, 85, 1, 4, 140, 0, 2, 
/* out0269_had-eta9-phi13*/	5, 84, 0, 2, 84, 1, 10, 84, 2, 1, 139, 0, 3, 140, 0, 1, 
/* out0270_had-eta10-phi13*/	4, 11, 0, 7, 28, 2, 2, 84, 1, 2, 139, 0, 5, 
/* out0271_had-eta11-phi13*/	2, 11, 0, 4, 11, 1, 5, 
/* out0272_had-eta12-phi13*/	4, 10, 0, 4, 11, 1, 4, 15, 8, 10, 15, 9, 1, 
/* out0273_had-eta13-phi13*/	4, 10, 0, 6, 10, 1, 10, 15, 8, 4, 15, 11, 3, 
/* out0274_had-eta14-phi13*/	3, 10, 1, 5, 10, 7, 13, 14, 9, 2, 
/* out0275_had-eta15-phi13*/	3, 10, 4, 3, 14, 8, 9, 14, 9, 5, 
/* out0276_had-eta16-phi13*/	3, 9, 0, 1, 14, 8, 7, 14, 11, 6, 
/* out0277_had-eta17-phi13*/	3, 9, 1, 5, 14, 5, 1, 14, 11, 5, 
/* out0278_had-eta18-phi13*/	3, 9, 7, 3, 12, 3, 1, 12, 5, 6, 
/* out0279_had-eta19-phi13*/	3, 12, 4, 2, 12, 5, 8, 12, 6, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 143, 0, 5, 
/* out0282_had-eta2-phi14*/	3, 88, 0, 3, 142, 0, 1, 143, 0, 3, 
/* out0283_had-eta3-phi14*/	4, 87, 0, 1, 88, 0, 8, 88, 1, 10, 142, 0, 5, 
/* out0284_had-eta4-phi14*/	6, 31, 0, 3, 31, 2, 4, 87, 0, 8, 87, 1, 7, 141, 0, 2, 142, 0, 2, 
/* out0285_had-eta5-phi14*/	7, 30, 0, 1, 31, 1, 4, 31, 2, 12, 86, 0, 7, 86, 1, 2, 87, 1, 1, 141, 0, 4, 
/* out0286_had-eta6-phi14*/	7, 30, 0, 3, 30, 1, 1, 30, 2, 14, 85, 0, 1, 86, 1, 4, 140, 0, 2, 141, 0, 2, 
/* out0287_had-eta7-phi14*/	7, 29, 0, 3, 29, 2, 3, 30, 1, 3, 30, 2, 2, 85, 0, 3, 85, 1, 3, 140, 0, 3, 
/* out0288_had-eta8-phi14*/	5, 29, 0, 1, 29, 1, 2, 29, 2, 12, 84, 0, 1, 140, 0, 2, 
/* out0289_had-eta9-phi14*/	8, 28, 0, 3, 28, 2, 4, 29, 1, 2, 29, 2, 1, 84, 0, 1, 84, 1, 1, 139, 0, 3, 140, 0, 1, 
/* out0290_had-eta10-phi14*/	3, 28, 1, 1, 28, 2, 9, 139, 0, 5, 
/* out0291_had-eta11-phi14*/	4, 15, 3, 9, 15, 9, 5, 28, 1, 3, 28, 2, 1, 
/* out0292_had-eta12-phi14*/	6, 15, 2, 4, 15, 3, 2, 15, 8, 2, 15, 9, 10, 15, 10, 11, 15, 11, 1, 
/* out0293_had-eta13-phi14*/	4, 15, 5, 6, 15, 6, 3, 15, 10, 5, 15, 11, 11, 
/* out0294_had-eta14-phi14*/	4, 14, 3, 10, 14, 9, 4, 15, 5, 6, 15, 11, 1, 
/* out0295_had-eta15-phi14*/	4, 14, 2, 3, 14, 3, 2, 14, 9, 5, 14, 10, 7, 
/* out0296_had-eta16-phi14*/	3, 14, 6, 4, 14, 10, 9, 14, 11, 3, 
/* out0297_had-eta17-phi14*/	2, 14, 5, 10, 14, 11, 2, 
/* out0298_had-eta18-phi14*/	2, 12, 3, 9, 14, 5, 1, 
/* out0299_had-eta19-phi14*/	4, 12, 2, 5, 12, 3, 2, 12, 5, 2, 12, 6, 15, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 148, 0, 5, 
/* out0302_had-eta2-phi15*/	4, 41, 0, 2, 41, 2, 1, 147, 0, 1, 148, 0, 3, 
/* out0303_had-eta3-phi15*/	5, 40, 0, 1, 41, 0, 1, 41, 1, 2, 41, 2, 15, 147, 0, 5, 
/* out0304_had-eta4-phi15*/	5, 31, 0, 8, 40, 0, 1, 40, 2, 14, 146, 0, 2, 147, 0, 2, 
/* out0305_had-eta5-phi15*/	8, 30, 0, 1, 31, 0, 5, 31, 1, 12, 39, 0, 1, 39, 2, 8, 40, 1, 1, 40, 2, 1, 146, 0, 4, 
/* out0306_had-eta6-phi15*/	6, 30, 0, 11, 30, 1, 6, 38, 2, 1, 39, 2, 4, 145, 0, 2, 146, 0, 2, 
/* out0307_had-eta7-phi15*/	4, 29, 0, 7, 30, 1, 6, 38, 2, 6, 145, 0, 3, 
/* out0308_had-eta8-phi15*/	4, 29, 0, 5, 29, 1, 9, 37, 2, 1, 145, 0, 2, 
/* out0309_had-eta9-phi15*/	5, 28, 0, 8, 29, 1, 3, 37, 2, 3, 144, 0, 3, 145, 0, 1, 
/* out0310_had-eta10-phi15*/	3, 28, 0, 4, 28, 1, 7, 144, 0, 5, 
/* out0311_had-eta11-phi15*/	4, 15, 0, 12, 15, 3, 3, 18, 2, 1, 28, 1, 4, 
/* out0312_had-eta12-phi15*/	6, 15, 0, 3, 15, 1, 8, 15, 2, 12, 15, 3, 2, 15, 6, 4, 15, 7, 1, 
/* out0313_had-eta13-phi15*/	4, 15, 4, 7, 15, 5, 3, 15, 6, 9, 15, 7, 5, 
/* out0314_had-eta14-phi15*/	4, 14, 0, 11, 14, 3, 3, 15, 4, 6, 15, 5, 1, 
/* out0315_had-eta15-phi15*/	4, 14, 0, 1, 14, 1, 3, 14, 2, 12, 14, 3, 1, 
/* out0316_had-eta16-phi15*/	3, 14, 2, 1, 14, 6, 12, 14, 7, 2, 
/* out0317_had-eta17-phi15*/	2, 14, 4, 8, 14, 5, 4, 
/* out0318_had-eta18-phi15*/	3, 12, 0, 6, 12, 3, 3, 14, 4, 1, 
/* out0319_had-eta19-phi15*/	4, 12, 0, 1, 12, 1, 1, 12, 2, 10, 12, 3, 1, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 148, 0, 5, 
/* out0322_had-eta2-phi16*/	3, 41, 0, 4, 147, 0, 1, 148, 0, 3, 
/* out0323_had-eta3-phi16*/	6, 40, 0, 2, 41, 0, 9, 41, 1, 14, 51, 0, 2, 51, 2, 10, 147, 0, 5, 
/* out0324_had-eta4-phi16*/	7, 40, 0, 12, 40, 1, 12, 40, 2, 1, 50, 2, 3, 51, 2, 4, 146, 0, 2, 147, 0, 2, 
/* out0325_had-eta5-phi16*/	6, 39, 0, 15, 39, 1, 4, 39, 2, 3, 40, 1, 3, 50, 2, 3, 146, 0, 4, 
/* out0326_had-eta6-phi16*/	7, 38, 0, 9, 38, 2, 1, 39, 1, 11, 39, 2, 1, 49, 2, 1, 145, 0, 2, 146, 0, 2, 
/* out0327_had-eta7-phi16*/	4, 38, 0, 4, 38, 1, 7, 38, 2, 7, 145, 0, 3, 
/* out0328_had-eta8-phi16*/	5, 37, 0, 7, 37, 2, 4, 38, 1, 3, 38, 2, 1, 145, 0, 2, 
/* out0329_had-eta9-phi16*/	5, 37, 0, 1, 37, 1, 4, 37, 2, 8, 144, 0, 3, 145, 0, 1, 
/* out0330_had-eta10-phi16*/	6, 18, 0, 3, 18, 2, 3, 28, 0, 1, 28, 1, 1, 37, 1, 2, 144, 0, 5, 
/* out0331_had-eta11-phi16*/	1, 18, 2, 9, 
/* out0332_had-eta12-phi16*/	7, 15, 0, 1, 15, 1, 8, 15, 7, 4, 16, 3, 2, 16, 9, 1, 18, 1, 1, 18, 2, 2, 
/* out0333_had-eta13-phi16*/	4, 15, 4, 3, 15, 7, 6, 16, 8, 4, 16, 9, 13, 
/* out0334_had-eta14-phi16*/	4, 14, 0, 3, 16, 8, 12, 16, 10, 1, 16, 11, 4, 
/* out0335_had-eta15-phi16*/	4, 14, 0, 1, 14, 1, 13, 14, 7, 1, 16, 11, 3, 
/* out0336_had-eta16-phi16*/	2, 13, 9, 1, 14, 7, 13, 
/* out0337_had-eta17-phi16*/	2, 13, 8, 5, 14, 4, 7, 
/* out0338_had-eta18-phi16*/	2, 12, 0, 7, 13, 8, 3, 
/* out0339_had-eta19-phi16*/	3, 12, 0, 2, 12, 1, 10, 12, 2, 1, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 153, 0, 5, 
/* out0342_had-eta2-phi17*/	2, 152, 0, 1, 153, 0, 3, 
/* out0343_had-eta3-phi17*/	7, 51, 0, 14, 51, 1, 8, 51, 2, 2, 60, 2, 2, 61, 0, 1, 61, 1, 16, 152, 0, 5, 
/* out0344_had-eta4-phi17*/	7, 50, 0, 15, 50, 1, 2, 50, 2, 4, 51, 1, 8, 60, 2, 5, 151, 0, 2, 152, 0, 2, 
/* out0345_had-eta5-phi17*/	6, 39, 1, 1, 49, 0, 7, 49, 2, 1, 50, 1, 12, 50, 2, 6, 151, 0, 4, 
/* out0346_had-eta6-phi17*/	6, 38, 0, 1, 49, 0, 3, 49, 1, 5, 49, 2, 13, 150, 0, 2, 151, 0, 2, 
/* out0347_had-eta7-phi17*/	7, 38, 0, 2, 38, 1, 5, 48, 0, 3, 48, 2, 7, 49, 1, 1, 49, 2, 1, 150, 0, 3, 
/* out0348_had-eta8-phi17*/	4, 37, 0, 7, 38, 1, 1, 48, 2, 7, 150, 0, 2, 
/* out0349_had-eta9-phi17*/	5, 37, 0, 1, 37, 1, 9, 47, 2, 3, 149, 0, 3, 150, 0, 1, 
/* out0350_had-eta10-phi17*/	4, 18, 0, 9, 37, 1, 1, 47, 2, 1, 149, 0, 5, 
/* out0351_had-eta11-phi17*/	3, 18, 0, 2, 18, 1, 6, 18, 2, 1, 
/* out0352_had-eta12-phi17*/	3, 16, 0, 5, 16, 3, 7, 18, 1, 4, 
/* out0353_had-eta13-phi17*/	4, 16, 2, 10, 16, 3, 7, 16, 9, 2, 16, 10, 6, 
/* out0354_had-eta14-phi17*/	4, 16, 5, 2, 16, 6, 6, 16, 10, 9, 16, 11, 4, 
/* out0355_had-eta15-phi17*/	3, 13, 3, 3, 16, 5, 9, 16, 11, 5, 
/* out0356_had-eta16-phi17*/	3, 13, 3, 4, 13, 9, 10, 13, 10, 1, 
/* out0357_had-eta17-phi17*/	3, 13, 8, 4, 13, 9, 5, 13, 10, 3, 
/* out0358_had-eta18-phi17*/	2, 13, 8, 4, 13, 11, 6, 
/* out0359_had-eta19-phi17*/	2, 12, 1, 5, 13, 11, 4, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 153, 0, 5, 
/* out0362_had-eta2-phi18*/	5, 61, 0, 2, 113, 0, 2, 113, 2, 1, 152, 0, 1, 153, 0, 3, 
/* out0363_had-eta3-phi18*/	6, 60, 0, 15, 60, 1, 1, 60, 2, 1, 61, 0, 13, 113, 2, 11, 152, 0, 5, 
/* out0364_had-eta4-phi18*/	9, 50, 0, 1, 50, 1, 1, 59, 0, 7, 59, 2, 1, 60, 0, 1, 60, 1, 15, 60, 2, 8, 151, 0, 2, 152, 0, 2, 
/* out0365_had-eta5-phi18*/	6, 49, 0, 3, 50, 1, 1, 59, 0, 3, 59, 1, 5, 59, 2, 15, 151, 0, 4, 
/* out0366_had-eta6-phi18*/	6, 49, 0, 3, 49, 1, 10, 58, 0, 2, 58, 2, 8, 150, 0, 2, 151, 0, 2, 
/* out0367_had-eta7-phi18*/	5, 48, 0, 13, 48, 1, 3, 48, 2, 1, 58, 2, 2, 150, 0, 3, 
/* out0368_had-eta8-phi18*/	4, 47, 0, 3, 48, 1, 11, 48, 2, 1, 150, 0, 2, 
/* out0369_had-eta9-phi18*/	5, 47, 0, 6, 47, 1, 1, 47, 2, 6, 149, 0, 3, 150, 0, 1, 
/* out0370_had-eta10-phi18*/	5, 17, 3, 2, 18, 0, 2, 47, 1, 3, 47, 2, 6, 149, 0, 5, 
/* out0371_had-eta11-phi18*/	4, 17, 3, 3, 17, 8, 3, 17, 9, 15, 18, 1, 4, 
/* out0372_had-eta12-phi18*/	4, 16, 0, 9, 17, 8, 13, 17, 11, 3, 18, 1, 1, 
/* out0373_had-eta13-phi18*/	5, 16, 0, 2, 16, 1, 13, 16, 2, 6, 16, 6, 2, 16, 7, 3, 
/* out0374_had-eta14-phi18*/	4, 16, 4, 5, 16, 5, 2, 16, 6, 8, 16, 7, 6, 
/* out0375_had-eta15-phi18*/	4, 13, 0, 5, 13, 3, 3, 16, 4, 6, 16, 5, 3, 
/* out0376_had-eta16-phi18*/	4, 13, 0, 1, 13, 2, 7, 13, 3, 6, 13, 10, 1, 
/* out0377_had-eta17-phi18*/	3, 13, 2, 3, 13, 6, 2, 13, 10, 8, 
/* out0378_had-eta18-phi18*/	4, 13, 5, 2, 13, 6, 2, 13, 10, 3, 13, 11, 3, 
/* out0379_had-eta19-phi18*/	2, 13, 5, 5, 13, 11, 3, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 158, 0, 5, 
/* out0382_had-eta2-phi19*/	3, 113, 0, 5, 157, 0, 1, 158, 0, 3, 
/* out0383_had-eta3-phi19*/	8, 111, 0, 9, 111, 2, 1, 112, 0, 1, 112, 2, 6, 113, 0, 9, 113, 1, 16, 113, 2, 4, 157, 0, 5, 
/* out0384_had-eta4-phi19*/	7, 59, 0, 4, 110, 0, 1, 111, 0, 5, 111, 1, 8, 111, 2, 15, 156, 0, 2, 157, 0, 2, 
/* out0385_had-eta5-phi19*/	6, 58, 0, 2, 59, 0, 2, 59, 1, 11, 110, 0, 2, 110, 2, 10, 156, 0, 4, 
/* out0386_had-eta6-phi19*/	6, 58, 0, 12, 58, 1, 7, 58, 2, 3, 110, 2, 1, 155, 0, 2, 156, 0, 2, 
/* out0387_had-eta7-phi19*/	6, 48, 1, 1, 57, 0, 6, 57, 2, 2, 58, 1, 6, 58, 2, 3, 155, 0, 3, 
/* out0388_had-eta8-phi19*/	4, 47, 0, 2, 48, 1, 1, 57, 2, 13, 155, 0, 2, 
/* out0389_had-eta9-phi19*/	5, 47, 0, 5, 47, 1, 6, 57, 2, 1, 154, 0, 3, 155, 0, 1, 
/* out0390_had-eta10-phi19*/	5, 17, 0, 11, 17, 3, 3, 47, 1, 6, 68, 2, 1, 154, 0, 5, 
/* out0391_had-eta11-phi19*/	7, 17, 0, 2, 17, 1, 1, 17, 2, 14, 17, 3, 8, 17, 6, 2, 17, 9, 1, 17, 10, 8, 
/* out0392_had-eta12-phi19*/	4, 17, 5, 6, 17, 6, 6, 17, 10, 8, 17, 11, 9, 
/* out0393_had-eta13-phi19*/	6, 16, 1, 3, 16, 7, 4, 17, 5, 4, 17, 11, 4, 19, 3, 3, 19, 9, 4, 
/* out0394_had-eta14-phi19*/	4, 16, 4, 4, 16, 7, 3, 19, 8, 6, 19, 9, 7, 
/* out0395_had-eta15-phi19*/	3, 13, 0, 8, 16, 4, 1, 19, 8, 7, 
/* out0396_had-eta16-phi19*/	3, 13, 0, 2, 13, 1, 8, 13, 2, 4, 
/* out0397_had-eta17-phi19*/	3, 13, 2, 2, 13, 6, 8, 13, 7, 2, 
/* out0398_had-eta18-phi19*/	3, 13, 4, 2, 13, 5, 4, 13, 6, 4, 
/* out0399_had-eta19-phi19*/	2, 13, 4, 2, 13, 5, 5, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 158, 0, 5, 
/* out0402_had-eta2-phi20*/	3, 112, 0, 6, 157, 0, 1, 158, 0, 3, 
/* out0403_had-eta3-phi20*/	6, 104, 0, 4, 111, 0, 1, 112, 0, 9, 112, 1, 16, 112, 2, 10, 157, 0, 5, 
/* out0404_had-eta4-phi20*/	7, 104, 0, 4, 104, 2, 15, 110, 0, 4, 111, 0, 1, 111, 1, 8, 156, 0, 2, 157, 0, 2, 
/* out0405_had-eta5-phi20*/	4, 110, 0, 9, 110, 1, 14, 110, 2, 4, 156, 0, 4, 
/* out0406_had-eta6-phi20*/	7, 58, 1, 2, 100, 0, 8, 100, 2, 8, 110, 1, 2, 110, 2, 1, 155, 0, 2, 156, 0, 2, 
/* out0407_had-eta7-phi20*/	5, 57, 0, 9, 57, 1, 1, 58, 1, 1, 100, 2, 8, 155, 0, 3, 
/* out0408_had-eta8-phi20*/	4, 57, 0, 1, 57, 1, 14, 68, 0, 1, 155, 0, 2, 
/* out0409_had-eta9-phi20*/	5, 57, 1, 1, 68, 0, 7, 68, 2, 5, 154, 0, 3, 155, 0, 1, 
/* out0410_had-eta10-phi20*/	4, 17, 0, 3, 17, 1, 1, 68, 2, 10, 154, 0, 5, 
/* out0411_had-eta11-phi20*/	4, 17, 1, 14, 17, 2, 2, 17, 6, 4, 17, 7, 13, 
/* out0412_had-eta12-phi20*/	5, 17, 4, 16, 17, 5, 5, 17, 6, 4, 17, 7, 3, 19, 0, 1, 
/* out0413_had-eta13-phi20*/	5, 17, 5, 1, 19, 0, 6, 19, 2, 4, 19, 3, 13, 19, 9, 1, 
/* out0414_had-eta14-phi20*/	4, 19, 2, 3, 19, 8, 1, 19, 9, 4, 19, 10, 13, 
/* out0415_had-eta15-phi20*/	3, 19, 8, 2, 19, 10, 2, 19, 11, 12, 
/* out0416_had-eta16-phi20*/	3, 13, 1, 8, 13, 7, 3, 19, 11, 3, 
/* out0417_had-eta17-phi20*/	2, 13, 4, 1, 13, 7, 11, 
/* out0418_had-eta18-phi20*/	1, 13, 4, 9, 
/* out0419_had-eta19-phi20*/	1, 13, 4, 2, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 163, 0, 5, 
/* out0422_had-eta2-phi21*/	3, 105, 0, 6, 162, 0, 1, 163, 0, 3, 
/* out0423_had-eta3-phi21*/	6, 102, 0, 1, 104, 0, 4, 105, 0, 9, 105, 1, 10, 105, 2, 16, 162, 0, 5, 
/* out0424_had-eta4-phi21*/	8, 101, 0, 4, 102, 0, 1, 102, 2, 8, 104, 0, 4, 104, 1, 16, 104, 2, 1, 161, 0, 2, 162, 0, 2, 
/* out0425_had-eta5-phi21*/	4, 101, 0, 9, 101, 1, 4, 101, 2, 14, 161, 0, 4, 
/* out0426_had-eta6-phi21*/	7, 70, 2, 2, 100, 0, 8, 100, 1, 8, 101, 1, 1, 101, 2, 2, 160, 0, 2, 161, 0, 2, 
/* out0427_had-eta7-phi21*/	5, 69, 0, 9, 69, 2, 1, 70, 2, 1, 100, 1, 8, 160, 0, 3, 
/* out0428_had-eta8-phi21*/	4, 68, 0, 1, 69, 0, 1, 69, 2, 14, 160, 0, 2, 
/* out0429_had-eta9-phi21*/	5, 68, 0, 7, 68, 1, 4, 69, 2, 1, 159, 0, 3, 160, 0, 1, 
/* out0430_had-eta10-phi21*/	4, 20, 0, 3, 20, 3, 1, 68, 1, 9, 159, 0, 5, 
/* out0431_had-eta11-phi21*/	5, 20, 2, 2, 20, 3, 14, 20, 9, 13, 20, 10, 4, 68, 1, 1, 
/* out0432_had-eta12-phi21*/	5, 19, 0, 2, 20, 8, 16, 20, 9, 3, 20, 10, 4, 20, 11, 5, 
/* out0433_had-eta13-phi21*/	4, 19, 0, 7, 19, 1, 12, 19, 2, 5, 20, 11, 1, 
/* out0434_had-eta14-phi21*/	4, 19, 2, 4, 19, 6, 13, 19, 7, 3, 19, 10, 1, 
/* out0435_had-eta15-phi21*/	4, 19, 4, 1, 19, 5, 13, 19, 6, 3, 19, 11, 1, 
/* out0436_had-eta16-phi21*/	3, 19, 5, 3, 21, 3, 8, 21, 9, 3, 
/* out0437_had-eta17-phi21*/	2, 21, 8, 1, 21, 9, 11, 
/* out0438_had-eta18-phi21*/	1, 21, 8, 9, 
/* out0439_had-eta19-phi21*/	1, 21, 8, 2, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 163, 0, 5, 
/* out0442_had-eta2-phi22*/	3, 103, 0, 5, 162, 0, 1, 163, 0, 3, 
/* out0443_had-eta3-phi22*/	8, 102, 0, 9, 102, 1, 1, 103, 0, 9, 103, 1, 4, 103, 2, 16, 105, 0, 1, 105, 1, 6, 162, 0, 5, 
/* out0444_had-eta4-phi22*/	7, 71, 0, 4, 101, 0, 1, 102, 0, 5, 102, 1, 15, 102, 2, 8, 161, 0, 2, 162, 0, 2, 
/* out0445_had-eta5-phi22*/	6, 70, 0, 2, 71, 0, 2, 71, 2, 11, 101, 0, 2, 101, 1, 10, 161, 0, 4, 
/* out0446_had-eta6-phi22*/	6, 70, 0, 12, 70, 1, 3, 70, 2, 7, 101, 1, 1, 160, 0, 2, 161, 0, 2, 
/* out0447_had-eta7-phi22*/	6, 69, 0, 6, 69, 1, 2, 70, 1, 3, 70, 2, 6, 80, 2, 1, 160, 0, 3, 
/* out0448_had-eta8-phi22*/	4, 69, 1, 13, 79, 0, 2, 80, 2, 1, 160, 0, 2, 
/* out0449_had-eta9-phi22*/	6, 68, 1, 1, 69, 1, 1, 79, 0, 5, 79, 2, 6, 159, 0, 3, 160, 0, 1, 
/* out0450_had-eta10-phi22*/	5, 20, 0, 11, 20, 1, 3, 68, 1, 1, 79, 2, 6, 159, 0, 5, 
/* out0451_had-eta11-phi22*/	7, 20, 0, 2, 20, 1, 8, 20, 2, 14, 20, 3, 1, 20, 6, 8, 20, 7, 1, 20, 10, 2, 
/* out0452_had-eta12-phi22*/	4, 20, 5, 9, 20, 6, 8, 20, 10, 6, 20, 11, 6, 
/* out0453_had-eta13-phi22*/	6, 19, 1, 4, 19, 7, 5, 20, 5, 4, 20, 11, 4, 22, 3, 3, 22, 9, 4, 
/* out0454_had-eta14-phi22*/	4, 19, 4, 6, 19, 7, 8, 22, 8, 4, 22, 9, 3, 
/* out0455_had-eta15-phi22*/	3, 19, 4, 9, 21, 0, 8, 22, 8, 1, 
/* out0456_had-eta16-phi22*/	3, 21, 0, 2, 21, 2, 4, 21, 3, 8, 
/* out0457_had-eta17-phi22*/	3, 21, 2, 2, 21, 9, 2, 21, 10, 8, 
/* out0458_had-eta18-phi22*/	3, 21, 8, 2, 21, 10, 4, 21, 11, 4, 
/* out0459_had-eta19-phi22*/	2, 21, 8, 2, 21, 11, 5, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 168, 0, 5, 
/* out0462_had-eta2-phi23*/	5, 73, 1, 2, 103, 0, 2, 103, 1, 1, 167, 0, 1, 168, 0, 3, 
/* out0463_had-eta3-phi23*/	6, 72, 0, 15, 72, 1, 1, 72, 2, 1, 73, 1, 13, 103, 1, 11, 167, 0, 5, 
/* out0464_had-eta4-phi23*/	9, 71, 0, 7, 71, 1, 1, 72, 0, 1, 72, 1, 8, 72, 2, 15, 82, 0, 1, 82, 2, 1, 166, 0, 2, 167, 0, 2, 
/* out0465_had-eta5-phi23*/	6, 71, 0, 3, 71, 1, 15, 71, 2, 5, 81, 0, 3, 82, 2, 1, 166, 0, 4, 
/* out0466_had-eta6-phi23*/	6, 70, 0, 2, 70, 1, 8, 81, 0, 3, 81, 2, 10, 165, 0, 2, 166, 0, 2, 
/* out0467_had-eta7-phi23*/	5, 70, 1, 2, 80, 0, 13, 80, 1, 1, 80, 2, 3, 165, 0, 3, 
/* out0468_had-eta8-phi23*/	4, 79, 0, 3, 80, 1, 1, 80, 2, 11, 165, 0, 2, 
/* out0469_had-eta9-phi23*/	5, 79, 0, 6, 79, 1, 6, 79, 2, 1, 164, 0, 3, 165, 0, 1, 
/* out0470_had-eta10-phi23*/	5, 20, 1, 2, 23, 0, 2, 79, 1, 6, 79, 2, 3, 164, 0, 5, 
/* out0471_had-eta11-phi23*/	4, 20, 1, 3, 20, 4, 3, 20, 7, 15, 23, 2, 4, 
/* out0472_had-eta12-phi23*/	4, 20, 4, 13, 20, 5, 3, 22, 0, 9, 23, 2, 1, 
/* out0473_had-eta13-phi23*/	5, 22, 0, 2, 22, 2, 6, 22, 3, 13, 22, 9, 3, 22, 10, 2, 
/* out0474_had-eta14-phi23*/	4, 22, 8, 5, 22, 9, 6, 22, 10, 8, 22, 11, 2, 
/* out0475_had-eta15-phi23*/	4, 21, 0, 5, 21, 1, 3, 22, 8, 6, 22, 11, 3, 
/* out0476_had-eta16-phi23*/	4, 21, 0, 1, 21, 1, 6, 21, 2, 7, 21, 6, 1, 
/* out0477_had-eta17-phi23*/	3, 21, 2, 3, 21, 6, 8, 21, 10, 2, 
/* out0478_had-eta18-phi23*/	4, 21, 5, 3, 21, 6, 3, 21, 10, 2, 21, 11, 2, 
/* out0479_had-eta19-phi23*/	2, 21, 5, 3, 21, 11, 5, 
/* out0480_had-eta0-phi24*/	0, 
/* out0481_had-eta1-phi24*/	1, 168, 0, 5, 
/* out0482_had-eta2-phi24*/	2, 167, 0, 1, 168, 0, 3, 
/* out0483_had-eta3-phi24*/	7, 72, 1, 2, 73, 0, 16, 73, 1, 1, 83, 0, 14, 83, 1, 2, 83, 2, 8, 167, 0, 5, 
/* out0484_had-eta4-phi24*/	7, 72, 1, 5, 82, 0, 15, 82, 1, 4, 82, 2, 2, 83, 2, 8, 166, 0, 2, 167, 0, 2, 
/* out0485_had-eta5-phi24*/	6, 81, 0, 7, 81, 1, 1, 82, 1, 6, 82, 2, 12, 91, 2, 1, 166, 0, 4, 
/* out0486_had-eta6-phi24*/	6, 81, 0, 3, 81, 1, 13, 81, 2, 5, 90, 0, 1, 165, 0, 2, 166, 0, 2, 
/* out0487_had-eta7-phi24*/	7, 80, 0, 3, 80, 1, 7, 81, 1, 1, 81, 2, 1, 90, 0, 2, 90, 2, 5, 165, 0, 3, 
/* out0488_had-eta8-phi24*/	4, 80, 1, 7, 89, 0, 7, 90, 2, 1, 165, 0, 2, 
/* out0489_had-eta9-phi24*/	5, 79, 1, 3, 89, 0, 1, 89, 2, 9, 164, 0, 3, 165, 0, 1, 
/* out0490_had-eta10-phi24*/	4, 23, 0, 9, 79, 1, 1, 89, 2, 1, 164, 0, 5, 
/* out0491_had-eta11-phi24*/	3, 23, 0, 2, 23, 1, 1, 23, 2, 6, 
/* out0492_had-eta12-phi24*/	3, 22, 0, 5, 22, 1, 7, 23, 2, 4, 
/* out0493_had-eta13-phi24*/	4, 22, 1, 7, 22, 2, 10, 22, 6, 6, 22, 7, 2, 
/* out0494_had-eta14-phi24*/	4, 22, 5, 4, 22, 6, 9, 22, 10, 6, 22, 11, 2, 
/* out0495_had-eta15-phi24*/	3, 21, 1, 3, 22, 5, 5, 22, 11, 9, 
/* out0496_had-eta16-phi24*/	3, 21, 1, 4, 21, 6, 1, 21, 7, 10, 
/* out0497_had-eta17-phi24*/	3, 21, 4, 4, 21, 6, 3, 21, 7, 5, 
/* out0498_had-eta18-phi24*/	2, 21, 4, 4, 21, 5, 6, 
/* out0499_had-eta19-phi24*/	1, 21, 5, 4, 
/* out0500_had-eta0-phi25*/	0, 
/* out0501_had-eta1-phi25*/	1, 173, 0, 5, 
/* out0502_had-eta2-phi25*/	3, 93, 0, 4, 172, 0, 1, 173, 0, 3, 
/* out0503_had-eta3-phi25*/	6, 83, 0, 2, 83, 1, 10, 92, 0, 2, 93, 0, 9, 93, 2, 14, 172, 0, 5, 
/* out0504_had-eta4-phi25*/	7, 82, 1, 3, 83, 1, 4, 92, 0, 12, 92, 1, 1, 92, 2, 12, 171, 0, 2, 172, 0, 2, 
/* out0505_had-eta5-phi25*/	6, 82, 1, 3, 91, 0, 15, 91, 1, 3, 91, 2, 4, 92, 2, 3, 171, 0, 4, 
/* out0506_had-eta6-phi25*/	7, 81, 1, 1, 90, 0, 9, 90, 1, 1, 91, 1, 1, 91, 2, 11, 170, 0, 2, 171, 0, 2, 
/* out0507_had-eta7-phi25*/	4, 90, 0, 4, 90, 1, 7, 90, 2, 7, 170, 0, 3, 
/* out0508_had-eta8-phi25*/	5, 89, 0, 7, 89, 1, 4, 90, 1, 1, 90, 2, 3, 170, 0, 2, 
/* out0509_had-eta9-phi25*/	5, 89, 0, 1, 89, 1, 8, 89, 2, 4, 169, 0, 3, 170, 0, 1, 
/* out0510_had-eta10-phi25*/	4, 23, 0, 3, 23, 1, 3, 89, 2, 2, 169, 0, 5, 
/* out0511_had-eta11-phi25*/	1, 23, 1, 9, 
/* out0512_had-eta12-phi25*/	4, 22, 1, 2, 22, 7, 1, 23, 1, 2, 23, 2, 1, 
/* out0513_had-eta13-phi25*/	2, 22, 4, 4, 22, 7, 13, 
/* out0514_had-eta14-phi25*/	3, 22, 4, 12, 22, 5, 4, 22, 6, 1, 
/* out0515_had-eta15-phi25*/	1, 22, 5, 3, 
/* out0516_had-eta16-phi25*/	1, 21, 7, 1, 
/* out0517_had-eta17-phi25*/	1, 21, 4, 5, 
/* out0518_had-eta18-phi25*/	1, 21, 4, 3, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	0, 
/* out0521_had-eta1-phi26*/	1, 173, 0, 5, 
/* out0522_had-eta2-phi26*/	4, 93, 0, 2, 93, 1, 1, 172, 0, 1, 173, 0, 3, 
/* out0523_had-eta3-phi26*/	5, 92, 0, 1, 93, 0, 1, 93, 1, 15, 93, 2, 2, 172, 0, 5, 
/* out0524_had-eta4-phi26*/	4, 92, 0, 1, 92, 1, 14, 171, 0, 2, 172, 0, 2, 
/* out0525_had-eta5-phi26*/	5, 91, 0, 1, 91, 1, 8, 92, 1, 1, 92, 2, 1, 171, 0, 4, 
/* out0526_had-eta6-phi26*/	4, 90, 1, 1, 91, 1, 4, 170, 0, 2, 171, 0, 2, 
/* out0527_had-eta7-phi26*/	2, 90, 1, 6, 170, 0, 3, 
/* out0528_had-eta8-phi26*/	2, 89, 1, 1, 170, 0, 2, 
/* out0529_had-eta9-phi26*/	3, 89, 1, 3, 169, 0, 3, 170, 0, 1, 
/* out0530_had-eta10-phi26*/	1, 169, 0, 5, 
/* out0531_had-eta11-phi26*/	1, 23, 1, 1, 
/* out0532_had-eta12-phi26*/	0, 
/* out0533_had-eta13-phi26*/	0, 
/* out0534_had-eta14-phi26*/	0, 
/* out0535_had-eta15-phi26*/	0, 
/* out0536_had-eta16-phi26*/	0, 
/* out0537_had-eta17-phi26*/	0, 
/* out0538_had-eta18-phi26*/	0, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	0, 
/* out0550_had-eta10-phi27*/	0, 
/* out0551_had-eta11-phi27*/	0, 
/* out0552_had-eta12-phi27*/	0, 
/* out0553_had-eta13-phi27*/	0, 
/* out0554_had-eta14-phi27*/	0, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	0, 
/* out0557_had-eta17-phi27*/	0, 
/* out0558_had-eta18-phi27*/	0, 
/* out0559_had-eta19-phi27*/	0, 
};