parameter integer matrixH [0:3902] = {
/* num inputs = 100(in0-in99) */
/* num outputs = 600(out0-out599) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1100 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	0,
/* out0006_em-eta6-phi0*/	0,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	0,
/* out0010_em-eta10-phi0*/	0,
/* out0011_em-eta11-phi0*/	0,
/* out0012_em-eta12-phi0*/	0,
/* out0013_em-eta13-phi0*/	0,
/* out0014_em-eta14-phi0*/	0,
/* out0015_em-eta15-phi0*/	0,
/* out0016_em-eta16-phi0*/	0,
/* out0017_em-eta17-phi0*/	0,
/* out0018_em-eta18-phi0*/	0,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	0,
/* out0026_em-eta6-phi1*/	0,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	0,
/* out0029_em-eta9-phi1*/	0,
/* out0030_em-eta10-phi1*/	0,
/* out0031_em-eta11-phi1*/	0,
/* out0032_em-eta12-phi1*/	0,
/* out0033_em-eta13-phi1*/	0,
/* out0034_em-eta14-phi1*/	0,
/* out0035_em-eta15-phi1*/	0,
/* out0036_em-eta16-phi1*/	0,
/* out0037_em-eta17-phi1*/	0,
/* out0038_em-eta18-phi1*/	0,
/* out0039_em-eta19-phi1*/	0,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	0,
/* out0046_em-eta6-phi2*/	0,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	0,
/* out0049_em-eta9-phi2*/	0,
/* out0050_em-eta10-phi2*/	0,
/* out0051_em-eta11-phi2*/	0,
/* out0052_em-eta12-phi2*/	0,
/* out0053_em-eta13-phi2*/	0,
/* out0054_em-eta14-phi2*/	0,
/* out0055_em-eta15-phi2*/	0,
/* out0056_em-eta16-phi2*/	0,
/* out0057_em-eta17-phi2*/	0,
/* out0058_em-eta18-phi2*/	0,
/* out0059_em-eta19-phi2*/	0,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	0,
/* out0065_em-eta5-phi3*/	2,79,0,4,79,2,4,
/* out0066_em-eta6-phi3*/	2,68,0,4,68,2,1,
/* out0067_em-eta7-phi3*/	2,57,0,1,68,2,3,
/* out0068_em-eta8-phi3*/	2,57,0,3,57,2,4,
/* out0069_em-eta9-phi3*/	1,46,0,2,
/* out0070_em-eta10-phi3*/	2,46,0,2,46,2,4,
/* out0071_em-eta11-phi3*/	1,35,0,1,
/* out0072_em-eta12-phi3*/	2,35,0,3,35,2,2,
/* out0073_em-eta13-phi3*/	1,35,2,2,
/* out0074_em-eta14-phi3*/	1,24,0,2,
/* out0075_em-eta15-phi3*/	2,24,0,2,24,2,2,
/* out0076_em-eta16-phi3*/	1,24,2,2,
/* out0077_em-eta17-phi3*/	1,14,2,1,
/* out0078_em-eta18-phi3*/	1,14,2,3,
/* out0079_em-eta19-phi3*/	1,14,0,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	3,79,0,3,79,1,1,89,2,2,
/* out0085_em-eta5-phi4*/	4,79,0,9,79,1,14,79,2,9,89,2,1,
/* out0086_em-eta6-phi4*/	6,68,0,12,68,1,9,68,2,2,79,2,3,80,0,1,80,2,1,
/* out0087_em-eta7-phi4*/	4,57,0,7,57,1,1,68,1,3,68,2,10,
/* out0088_em-eta8-phi4*/	3,57,0,5,57,1,6,57,2,7,
/* out0089_em-eta9-phi4*/	3,46,0,9,46,1,1,57,2,5,
/* out0090_em-eta10-phi4*/	3,46,0,3,46,1,3,46,2,7,
/* out0091_em-eta11-phi4*/	2,35,0,7,46,2,4,
/* out0092_em-eta12-phi4*/	3,35,0,4,35,1,1,35,2,4,
/* out0093_em-eta13-phi4*/	2,24,0,1,35,2,6,
/* out0094_em-eta14-phi4*/	1,24,0,6,
/* out0095_em-eta15-phi4*/	2,24,0,2,24,2,3,
/* out0096_em-eta16-phi4*/	1,24,2,4,
/* out0097_em-eta17-phi4*/	2,14,2,4,24,2,1,
/* out0098_em-eta18-phi4*/	2,14,0,1,14,2,3,
/* out0099_em-eta19-phi4*/	1,14,0,1,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	2,89,1,3,89,2,8,
/* out0105_em-eta5-phi5*/	5,79,1,1,80,0,14,80,1,4,89,1,11,89,2,5,
/* out0106_em-eta6-phi5*/	5,68,1,3,69,0,5,80,0,1,80,1,2,80,2,15,
/* out0107_em-eta7-phi5*/	5,57,1,1,68,1,1,69,0,10,69,1,1,69,2,9,
/* out0108_em-eta8-phi5*/	3,57,1,7,58,0,8,69,2,4,
/* out0109_em-eta9-phi5*/	4,46,1,4,57,1,1,58,0,3,58,2,8,
/* out0110_em-eta10-phi5*/	3,46,1,8,47,0,4,58,2,1,
/* out0111_em-eta11-phi5*/	5,35,0,1,35,1,3,46,2,1,47,0,2,47,2,3,
/* out0112_em-eta12-phi5*/	1,35,1,9,
/* out0113_em-eta13-phi5*/	5,24,0,1,35,1,2,35,2,2,36,0,1,36,2,1,
/* out0114_em-eta14-phi5*/	2,24,0,2,24,1,4,
/* out0115_em-eta15-phi5*/	2,24,1,5,24,2,1,
/* out0116_em-eta16-phi5*/	2,24,1,1,24,2,3,
/* out0117_em-eta17-phi5*/	2,14,0,1,14,2,4,
/* out0118_em-eta18-phi5*/	2,14,0,3,14,2,1,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	3,89,1,2,90,0,5,90,1,4,
/* out0125_em-eta5-phi6*/	5,80,1,5,81,0,3,90,0,11,90,1,5,90,2,15,
/* out0126_em-eta6-phi6*/	5,69,0,1,69,1,2,80,1,5,81,0,11,81,2,8,
/* out0127_em-eta7-phi6*/	4,69,1,13,69,2,1,70,0,5,81,2,2,
/* out0128_em-eta8-phi6*/	5,58,0,5,58,1,7,69,2,2,70,0,1,70,2,3,
/* out0129_em-eta9-phi6*/	2,58,1,7,58,2,7,
/* out0130_em-eta10-phi6*/	2,47,0,9,47,1,3,
/* out0131_em-eta11-phi6*/	3,47,0,1,47,1,1,47,2,9,
/* out0132_em-eta12-phi6*/	3,35,1,1,36,0,6,47,2,2,
/* out0133_em-eta13-phi6*/	2,36,0,4,36,2,3,
/* out0134_em-eta14-phi6*/	2,24,1,2,36,2,4,
/* out0135_em-eta15-phi6*/	2,24,1,3,25,0,2,
/* out0136_em-eta16-phi6*/	2,24,1,1,25,0,2,
/* out0137_em-eta17-phi6*/	2,14,0,3,25,2,1,
/* out0138_em-eta18-phi6*/	1,14,0,4,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	2,90,1,1,91,0,2,
/* out0145_em-eta5-phi7*/	6,81,0,1,81,1,2,90,1,6,90,2,1,91,0,13,91,2,8,
/* out0146_em-eta6-phi7*/	5,81,0,1,81,1,14,81,2,4,82,0,5,91,2,2,
/* out0147_em-eta7-phi7*/	4,70,0,10,70,1,8,81,2,2,82,2,1,
/* out0148_em-eta8-phi7*/	4,58,1,1,59,0,3,70,1,2,70,2,12,
/* out0149_em-eta9-phi7*/	3,58,1,1,59,0,11,59,2,4,
/* out0150_em-eta10-phi7*/	3,47,1,6,48,0,1,59,2,5,
/* out0151_em-eta11-phi7*/	3,47,1,6,47,2,2,48,0,3,
/* out0152_em-eta12-phi7*/	3,36,0,4,36,1,4,48,2,1,
/* out0153_em-eta13-phi7*/	3,36,0,1,36,1,4,36,2,2,
/* out0154_em-eta14-phi7*/	2,25,0,1,36,2,5,
/* out0155_em-eta15-phi7*/	1,25,0,5,
/* out0156_em-eta16-phi7*/	2,25,0,3,25,2,2,
/* out0157_em-eta17-phi7*/	1,25,2,3,
/* out0158_em-eta18-phi7*/	2,14,0,2,25,2,1,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	5,91,0,1,91,1,1,97,0,11,97,1,5,97,2,8,
/* out0165_em-eta5-phi8*/	7,91,1,15,91,2,5,92,0,8,92,2,2,97,0,4,97,1,8,97,2,4,
/* out0166_em-eta6-phi8*/	5,82,0,11,82,1,11,82,2,3,91,2,1,92,2,1,
/* out0167_em-eta7-phi8*/	3,70,1,4,71,0,7,82,2,11,
/* out0168_em-eta8-phi8*/	6,59,0,1,59,1,3,70,1,2,70,2,1,71,0,5,71,2,6,
/* out0169_em-eta9-phi8*/	3,59,0,1,59,1,12,59,2,2,
/* out0170_em-eta10-phi8*/	4,48,0,6,48,1,1,59,1,1,59,2,5,
/* out0171_em-eta11-phi8*/	3,48,0,6,48,1,1,48,2,4,
/* out0172_em-eta12-phi8*/	2,36,1,2,48,2,6,
/* out0173_em-eta13-phi8*/	2,36,1,5,37,0,3,
/* out0174_em-eta14-phi8*/	6,25,0,1,25,1,1,36,1,1,36,2,1,37,0,1,37,2,1,
/* out0175_em-eta15-phi8*/	2,25,0,2,25,1,4,
/* out0176_em-eta16-phi8*/	2,25,1,2,25,2,2,
/* out0177_em-eta17-phi8*/	1,25,2,4,
/* out0178_em-eta18-phi8*/	1,25,2,1,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	6,97,0,1,97,1,2,97,2,3,98,0,5,98,1,1,98,2,3,
/* out0185_em-eta5-phi9*/	8,92,0,8,92,1,16,92,2,6,97,1,1,97,2,1,98,0,7,98,1,7,98,2,1,
/* out0186_em-eta6-phi9*/	4,82,1,4,83,0,15,83,2,1,92,2,7,
/* out0187_em-eta7-phi9*/	6,71,0,3,71,1,9,82,1,1,82,2,1,83,0,1,83,2,7,
/* out0188_em-eta8-phi9*/	4,60,0,2,71,0,1,71,1,7,71,2,9,
/* out0189_em-eta9-phi9*/	3,60,0,13,60,2,1,71,2,1,
/* out0190_em-eta10-phi9*/	3,48,1,5,60,0,1,60,2,7,
/* out0191_em-eta11-phi9*/	2,48,1,9,48,2,1,
/* out0192_em-eta12-phi9*/	2,37,0,4,48,2,4,
/* out0193_em-eta13-phi9*/	1,37,0,7,
/* out0194_em-eta14-phi9*/	2,37,0,1,37,2,6,
/* out0195_em-eta15-phi9*/	2,25,1,4,37,2,1,
/* out0196_em-eta16-phi9*/	1,25,1,4,
/* out0197_em-eta17-phi9*/	2,25,1,1,25,2,2,
/* out0198_em-eta18-phi9*/	0,
/* out0199_em-eta19-phi9*/	0,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	6,98,0,3,98,1,1,98,2,5,99,0,3,99,1,2,99,2,1,
/* out0205_em-eta5-phi10*/	8,93,0,16,93,1,8,93,2,6,98,0,1,98,1,7,98,2,7,99,0,1,99,1,1,
/* out0206_em-eta6-phi10*/	4,83,1,15,83,2,1,84,0,4,93,2,7,
/* out0207_em-eta7-phi10*/	6,72,0,9,72,1,3,83,1,1,83,2,7,84,0,1,84,2,1,
/* out0208_em-eta8-phi10*/	4,60,1,2,72,0,7,72,1,1,72,2,9,
/* out0209_em-eta9-phi10*/	3,60,1,13,60,2,1,72,2,1,
/* out0210_em-eta10-phi10*/	3,49,0,5,60,1,1,60,2,7,
/* out0211_em-eta11-phi10*/	2,49,0,9,49,2,1,
/* out0212_em-eta12-phi10*/	2,37,1,4,49,2,4,
/* out0213_em-eta13-phi10*/	1,37,1,7,
/* out0214_em-eta14-phi10*/	2,37,1,1,37,2,6,
/* out0215_em-eta15-phi10*/	2,26,0,4,37,2,1,
/* out0216_em-eta16-phi10*/	1,26,0,4,
/* out0217_em-eta17-phi10*/	2,26,0,1,26,2,2,
/* out0218_em-eta18-phi10*/	0,
/* out0219_em-eta19-phi10*/	0,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	5,94,0,1,94,1,1,99,0,8,99,1,5,99,2,11,
/* out0225_em-eta5-phi11*/	7,93,1,8,93,2,2,94,0,15,94,2,5,99,0,4,99,1,8,99,2,4,
/* out0226_em-eta6-phi11*/	5,84,0,11,84,1,11,84,2,3,93,2,1,94,2,1,
/* out0227_em-eta7-phi11*/	3,72,1,7,73,0,4,84,2,11,
/* out0228_em-eta8-phi11*/	6,61,0,3,61,1,1,72,1,5,72,2,6,73,0,2,73,2,1,
/* out0229_em-eta9-phi11*/	3,61,0,12,61,1,1,61,2,2,
/* out0230_em-eta10-phi11*/	4,49,0,1,49,1,6,61,0,1,61,2,5,
/* out0231_em-eta11-phi11*/	3,49,0,1,49,1,6,49,2,4,
/* out0232_em-eta12-phi11*/	2,38,0,2,49,2,6,
/* out0233_em-eta13-phi11*/	2,37,1,3,38,0,5,
/* out0234_em-eta14-phi11*/	6,26,0,1,26,1,1,37,1,1,37,2,1,38,0,1,38,2,1,
/* out0235_em-eta15-phi11*/	2,26,0,4,26,1,2,
/* out0236_em-eta16-phi11*/	2,26,0,2,26,2,2,
/* out0237_em-eta17-phi11*/	1,26,2,4,
/* out0238_em-eta18-phi11*/	1,26,2,1,
/* out0239_em-eta19-phi11*/	0,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	2,94,1,2,95,1,1,
/* out0245_em-eta5-phi12*/	7,85,0,2,85,1,1,94,1,13,94,2,8,95,0,13,95,1,1,95,2,1,
/* out0246_em-eta6-phi12*/	5,84,1,5,85,0,14,85,1,1,85,2,4,94,2,2,
/* out0247_em-eta7-phi12*/	4,73,0,8,73,1,10,84,2,1,85,2,2,
/* out0248_em-eta8-phi12*/	4,61,1,3,62,0,1,73,0,2,73,2,12,
/* out0249_em-eta9-phi12*/	3,61,1,11,61,2,4,62,0,1,
/* out0250_em-eta10-phi12*/	3,49,1,1,50,0,6,61,2,5,
/* out0251_em-eta11-phi12*/	3,49,1,3,50,0,6,50,2,2,
/* out0252_em-eta12-phi12*/	3,38,0,4,38,1,4,49,2,1,
/* out0253_em-eta13-phi12*/	3,38,0,4,38,1,1,38,2,2,
/* out0254_em-eta14-phi12*/	2,26,1,1,38,2,5,
/* out0255_em-eta15-phi12*/	1,26,1,5,
/* out0256_em-eta16-phi12*/	2,26,1,3,26,2,2,
/* out0257_em-eta17-phi12*/	1,26,2,3,
/* out0258_em-eta18-phi12*/	2,15,1,2,26,2,1,
/* out0259_em-eta19-phi12*/	0,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	2,95,1,6,96,0,2,
/* out0265_em-eta5-phi13*/	5,85,1,3,86,0,5,95,0,3,95,1,8,95,2,15,
/* out0266_em-eta6-phi13*/	5,74,0,2,74,1,1,85,1,11,85,2,8,86,0,5,
/* out0267_em-eta7-phi13*/	4,73,1,5,74,0,13,74,2,1,85,2,2,
/* out0268_em-eta8-phi13*/	5,62,0,7,62,1,5,73,1,1,73,2,3,74,2,2,
/* out0269_em-eta9-phi13*/	2,62,0,7,62,2,7,
/* out0270_em-eta10-phi13*/	2,50,0,3,50,1,9,
/* out0271_em-eta11-phi13*/	3,50,0,1,50,1,1,50,2,9,
/* out0272_em-eta12-phi13*/	3,38,1,6,39,0,1,50,2,2,
/* out0273_em-eta13-phi13*/	2,38,1,4,38,2,3,
/* out0274_em-eta14-phi13*/	2,27,0,2,38,2,4,
/* out0275_em-eta15-phi13*/	2,26,1,2,27,0,3,
/* out0276_em-eta16-phi13*/	2,26,1,2,27,0,1,
/* out0277_em-eta17-phi13*/	2,15,1,3,26,2,1,
/* out0278_em-eta18-phi13*/	1,15,1,4,
/* out0279_em-eta19-phi13*/	0,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	2,96,0,10,96,2,1,
/* out0285_em-eta5-phi14*/	5,86,0,4,86,1,14,87,0,1,96,0,4,96,2,13,
/* out0286_em-eta6-phi14*/	5,74,1,5,75,0,3,86,0,2,86,1,1,86,2,15,
/* out0287_em-eta7-phi14*/	5,63,0,1,74,0,1,74,1,10,74,2,9,75,0,1,
/* out0288_em-eta8-phi14*/	3,62,1,8,63,0,7,74,2,4,
/* out0289_em-eta9-phi14*/	4,51,0,4,62,1,3,62,2,8,63,0,1,
/* out0290_em-eta10-phi14*/	3,50,1,4,51,0,8,62,2,1,
/* out0291_em-eta11-phi14*/	5,39,0,3,39,1,1,50,1,2,50,2,3,51,2,1,
/* out0292_em-eta12-phi14*/	1,39,0,9,
/* out0293_em-eta13-phi14*/	5,27,1,1,38,1,1,38,2,1,39,0,2,39,2,2,
/* out0294_em-eta14-phi14*/	2,27,0,4,27,1,2,
/* out0295_em-eta15-phi14*/	2,27,0,5,27,2,1,
/* out0296_em-eta16-phi14*/	2,27,0,1,27,2,3,
/* out0297_em-eta17-phi14*/	2,15,1,1,15,2,4,
/* out0298_em-eta18-phi14*/	2,15,1,3,15,2,1,
/* out0299_em-eta19-phi14*/	0,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	3,87,0,1,87,1,3,96,2,1,
/* out0305_em-eta5-phi15*/	4,87,0,14,87,1,9,87,2,9,96,2,1,
/* out0306_em-eta6-phi15*/	6,75,0,9,75,1,12,75,2,2,86,1,1,86,2,1,87,2,3,
/* out0307_em-eta7-phi15*/	4,63,0,1,63,1,7,75,0,3,75,2,10,
/* out0308_em-eta8-phi15*/	3,63,0,6,63,1,5,63,2,7,
/* out0309_em-eta9-phi15*/	3,51,0,1,51,1,9,63,2,5,
/* out0310_em-eta10-phi15*/	3,51,0,3,51,1,3,51,2,7,
/* out0311_em-eta11-phi15*/	2,39,1,7,51,2,4,
/* out0312_em-eta12-phi15*/	3,39,0,1,39,1,4,39,2,4,
/* out0313_em-eta13-phi15*/	2,27,1,1,39,2,6,
/* out0314_em-eta14-phi15*/	1,27,1,6,
/* out0315_em-eta15-phi15*/	2,27,1,2,27,2,3,
/* out0316_em-eta16-phi15*/	1,27,2,4,
/* out0317_em-eta17-phi15*/	2,15,2,4,27,2,1,
/* out0318_em-eta18-phi15*/	2,15,1,1,15,2,3,
/* out0319_em-eta19-phi15*/	1,15,1,1,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	1,88,0,7,
/* out0325_em-eta5-phi16*/	6,76,0,5,76,1,7,87,1,4,87,2,4,88,0,8,88,2,8,
/* out0326_em-eta6-phi16*/	6,64,1,2,75,1,4,75,2,1,76,0,11,76,1,1,76,2,7,
/* out0327_em-eta7-phi16*/	5,63,1,1,64,0,14,64,1,4,64,2,1,75,2,3,
/* out0328_em-eta8-phi16*/	6,52,0,4,52,1,3,63,1,3,63,2,4,64,0,2,64,2,3,
/* out0329_em-eta9-phi16*/	3,51,1,2,52,0,11,52,2,1,
/* out0330_em-eta10-phi16*/	6,40,0,4,40,1,1,51,1,2,51,2,4,52,0,1,52,2,1,
/* out0331_em-eta11-phi16*/	2,39,1,1,40,0,9,
/* out0332_em-eta12-phi16*/	5,28,0,1,39,1,3,39,2,2,40,0,1,40,2,1,
/* out0333_em-eta13-phi16*/	2,28,0,6,39,2,2,
/* out0334_em-eta14-phi16*/	2,27,1,2,28,0,4,
/* out0335_em-eta15-phi16*/	3,16,0,1,27,1,2,27,2,2,
/* out0336_em-eta16-phi16*/	2,16,0,3,27,2,2,
/* out0337_em-eta17-phi16*/	2,15,2,1,16,0,3,
/* out0338_em-eta18-phi16*/	1,15,2,3,
/* out0339_em-eta19-phi16*/	1,15,1,1,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	4,77,0,1,77,1,4,88,0,1,88,2,3,
/* out0345_em-eta5-phi17*/	5,76,1,7,77,0,15,77,1,3,77,2,4,88,2,5,
/* out0346_em-eta6-phi17*/	5,64,1,2,65,0,12,65,1,2,76,1,1,76,2,9,
/* out0347_em-eta7-phi17*/	4,53,0,3,64,1,8,64,2,8,65,0,3,
/* out0348_em-eta8-phi17*/	3,52,1,9,53,0,5,64,2,4,
/* out0349_em-eta9-phi17*/	2,52,1,4,52,2,11,
/* out0350_em-eta10-phi17*/	3,40,1,10,41,0,1,52,2,2,
/* out0351_em-eta11-phi17*/	3,40,0,2,40,1,2,40,2,6,
/* out0352_em-eta12-phi17*/	2,28,1,5,40,2,4,
/* out0353_em-eta13-phi17*/	3,28,0,3,28,1,4,28,2,1,
/* out0354_em-eta14-phi17*/	2,28,0,2,28,2,4,
/* out0355_em-eta15-phi17*/	3,16,0,1,16,1,3,28,2,1,
/* out0356_em-eta16-phi17*/	2,16,0,3,16,1,1,
/* out0357_em-eta17-phi17*/	1,16,0,3,
/* out0358_em-eta18-phi17*/	2,16,0,2,16,2,1,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	4,77,1,4,78,0,12,78,1,6,78,2,7,
/* out0365_em-eta5-phi18*/	8,65,1,1,66,0,10,66,1,2,77,1,5,77,2,12,78,0,2,78,1,7,78,2,5,
/* out0366_em-eta6-phi18*/	5,54,0,1,65,0,1,65,1,13,65,2,9,66,0,3,
/* out0367_em-eta7-phi18*/	4,53,0,1,53,1,12,54,0,2,65,2,7,
/* out0368_em-eta8-phi18*/	3,53,0,7,53,1,1,53,2,10,
/* out0369_em-eta9-phi18*/	4,41,0,7,41,1,7,52,2,1,53,2,1,
/* out0370_em-eta10-phi18*/	3,40,1,2,41,0,8,41,2,3,
/* out0371_em-eta11-phi18*/	4,29,0,4,29,1,1,40,1,1,40,2,4,
/* out0372_em-eta12-phi18*/	3,28,1,3,29,0,5,40,2,1,
/* out0373_em-eta13-phi18*/	2,28,1,4,28,2,3,
/* out0374_em-eta14-phi18*/	1,28,2,6,
/* out0375_em-eta15-phi18*/	2,16,1,4,28,2,1,
/* out0376_em-eta16-phi18*/	2,16,1,4,16,2,1,
/* out0377_em-eta17-phi18*/	1,16,2,3,
/* out0378_em-eta18-phi18*/	1,16,2,3,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	3,67,1,9,78,0,2,78,2,2,
/* out0385_em-eta5-phi19*/	9,55,0,1,66,0,2,66,1,14,66,2,9,67,0,16,67,1,1,67,2,1,78,1,3,78,2,2,
/* out0386_em-eta6-phi19*/	5,54,0,4,54,1,13,55,0,1,66,0,1,66,2,7,
/* out0387_em-eta7-phi19*/	4,42,1,2,53,1,3,54,0,9,54,2,8,
/* out0388_em-eta8-phi19*/	3,42,0,10,42,1,2,53,2,5,
/* out0389_em-eta9-phi19*/	3,41,1,9,41,2,3,42,0,3,
/* out0390_em-eta10-phi19*/	3,29,1,2,30,0,1,41,2,10,
/* out0391_em-eta11-phi19*/	2,29,0,2,29,1,9,
/* out0392_em-eta12-phi19*/	2,29,0,4,29,2,5,
/* out0393_em-eta13-phi19*/	4,17,0,2,17,1,3,29,0,1,29,2,2,
/* out0394_em-eta14-phi19*/	1,17,0,6,
/* out0395_em-eta15-phi19*/	2,16,1,1,17,0,4,
/* out0396_em-eta16-phi19*/	2,16,1,3,16,2,2,
/* out0397_em-eta17-phi19*/	1,16,2,4,
/* out0398_em-eta18-phi19*/	1,16,2,2,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	3,56,1,2,67,1,6,67,2,2,
/* out0405_em-eta5-phi20*/	6,55,0,5,55,1,14,55,2,2,56,0,5,56,1,4,67,2,13,
/* out0406_em-eta6-phi20*/	6,43,0,1,43,1,4,54,1,3,54,2,2,55,0,9,55,2,8,
/* out0407_em-eta7-phi20*/	3,42,1,4,43,0,11,54,2,6,
/* out0408_em-eta8-phi20*/	3,42,0,2,42,1,8,42,2,9,
/* out0409_em-eta9-phi20*/	4,30,0,2,30,1,7,42,0,1,42,2,6,
/* out0410_em-eta10-phi20*/	3,30,0,11,30,1,1,30,2,1,
/* out0411_em-eta11-phi20*/	5,18,0,1,29,1,4,29,2,3,30,0,2,30,2,1,
/* out0412_em-eta12-phi20*/	2,18,0,2,29,2,6,
/* out0413_em-eta13-phi20*/	1,17,1,7,
/* out0414_em-eta14-phi20*/	3,17,0,2,17,1,2,17,2,2,
/* out0415_em-eta15-phi20*/	2,17,0,2,17,2,3,
/* out0416_em-eta16-phi20*/	3,7,1,1,7,2,1,17,2,1,
/* out0417_em-eta17-phi20*/	1,7,1,3,
/* out0418_em-eta18-phi20*/	1,7,1,2,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	1,56,1,4,
/* out0425_em-eta5-phi21*/	7,44,0,4,44,1,8,55,1,2,55,2,3,56,0,11,56,1,6,56,2,16,
/* out0426_em-eta6-phi21*/	4,43,1,10,43,2,1,44,0,12,55,2,3,
/* out0427_em-eta7-phi21*/	4,31,1,1,43,0,3,43,1,2,43,2,15,
/* out0428_em-eta8-phi21*/	4,31,0,9,31,1,7,42,2,1,43,0,1,
/* out0429_em-eta9-phi21*/	3,30,1,7,30,2,1,31,0,7,
/* out0430_em-eta10-phi21*/	2,30,1,1,30,2,11,
/* out0431_em-eta11-phi21*/	3,18,0,1,18,1,7,30,2,2,
/* out0432_em-eta12-phi21*/	2,18,0,8,18,1,1,
/* out0433_em-eta13-phi21*/	2,17,1,4,18,0,4,
/* out0434_em-eta14-phi21*/	1,17,2,6,
/* out0435_em-eta15-phi21*/	2,7,2,1,17,2,4,
/* out0436_em-eta16-phi21*/	1,7,2,5,
/* out0437_em-eta17-phi21*/	1,7,1,3,
/* out0438_em-eta18-phi21*/	1,7,1,2,
/* out0439_em-eta19-phi21*/	0,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	1,45,1,5,
/* out0445_em-eta5-phi22*/	7,33,0,3,33,1,2,44,1,8,44,2,4,45,0,16,45,1,10,45,2,9,
/* out0446_em-eta6-phi22*/	4,32,0,1,32,1,10,33,0,3,44,2,12,
/* out0447_em-eta7-phi22*/	4,31,1,1,32,0,15,32,1,2,32,2,3,
/* out0448_em-eta8-phi22*/	4,20,0,1,31,1,7,31,2,9,32,2,1,
/* out0449_em-eta9-phi22*/	3,19,0,1,19,1,7,31,2,7,
/* out0450_em-eta10-phi22*/	2,19,0,11,19,1,1,
/* out0451_em-eta11-phi22*/	3,18,1,7,18,2,1,19,0,2,
/* out0452_em-eta12-phi22*/	2,18,1,1,18,2,8,
/* out0453_em-eta13-phi22*/	2,8,1,4,18,2,4,
/* out0454_em-eta14-phi22*/	1,8,0,6,
/* out0455_em-eta15-phi22*/	2,7,2,1,8,0,4,
/* out0456_em-eta16-phi22*/	1,7,2,5,
/* out0457_em-eta17-phi22*/	3,7,0,3,7,1,2,7,2,1,
/* out0458_em-eta18-phi22*/	1,7,1,2,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	3,34,1,8,45,1,1,45,2,1,
/* out0465_em-eta5-phi23*/	7,33,0,2,33,1,14,33,2,5,34,0,16,34,1,5,34,2,2,45,2,6,
/* out0466_em-eta6-phi23*/	6,21,0,2,21,1,3,32,1,4,32,2,1,33,0,8,33,2,9,
/* out0467_em-eta7-phi23*/	3,20,1,4,21,0,6,32,2,11,
/* out0468_em-eta8-phi23*/	3,20,0,9,20,1,8,20,2,2,
/* out0469_em-eta9-phi23*/	4,19,1,7,19,2,2,20,0,6,20,2,1,
/* out0470_em-eta10-phi23*/	3,19,0,1,19,1,1,19,2,11,
/* out0471_em-eta11-phi23*/	5,9,0,3,9,1,4,18,2,1,19,0,1,19,2,2,
/* out0472_em-eta12-phi23*/	2,9,0,6,18,2,2,
/* out0473_em-eta13-phi23*/	1,8,1,7,
/* out0474_em-eta14-phi23*/	3,8,0,2,8,1,2,8,2,2,
/* out0475_em-eta15-phi23*/	2,8,0,3,8,2,2,
/* out0476_em-eta16-phi23*/	3,7,0,3,7,2,2,8,0,1,
/* out0477_em-eta17-phi23*/	1,7,0,8,
/* out0478_em-eta18-phi23*/	2,7,0,1,7,1,1,
/* out0479_em-eta19-phi23*/	0,
/* out0480_em-eta0-phi24*/	0,
/* out0481_em-eta1-phi24*/	0,
/* out0482_em-eta2-phi24*/	0,
/* out0483_em-eta3-phi24*/	0,
/* out0484_em-eta4-phi24*/	4,23,0,2,23,2,2,34,1,3,34,2,6,
/* out0485_em-eta5-phi24*/	7,22,0,9,22,1,14,22,2,2,23,0,2,23,1,3,33,2,1,34,2,8,
/* out0486_em-eta6-phi24*/	5,21,1,13,21,2,4,22,0,7,22,2,1,33,2,1,
/* out0487_em-eta7-phi24*/	4,11,1,3,20,1,2,21,0,8,21,2,9,
/* out0488_em-eta8-phi24*/	3,11,0,5,20,1,2,20,2,10,
/* out0489_em-eta9-phi24*/	3,10,0,3,10,1,9,20,2,3,
/* out0490_em-eta10-phi24*/	3,9,1,2,10,0,10,19,2,1,
/* out0491_em-eta11-phi24*/	2,9,1,9,9,2,2,
/* out0492_em-eta12-phi24*/	2,9,0,5,9,2,4,
/* out0493_em-eta13-phi24*/	4,8,1,3,8,2,2,9,0,2,9,2,1,
/* out0494_em-eta14-phi24*/	1,8,2,6,
/* out0495_em-eta15-phi24*/	2,0,1,1,8,2,4,
/* out0496_em-eta16-phi24*/	2,0,0,2,0,1,3,
/* out0497_em-eta17-phi24*/	1,0,0,4,
/* out0498_em-eta18-phi24*/	2,0,0,2,7,0,1,
/* out0499_em-eta19-phi24*/	0,
/* out0500_em-eta0-phi25*/	0,
/* out0501_em-eta1-phi25*/	0,
/* out0502_em-eta2-phi25*/	0,
/* out0503_em-eta3-phi25*/	0,
/* out0504_em-eta4-phi25*/	4,13,1,4,23,0,7,23,1,6,23,2,12,
/* out0505_em-eta5-phi25*/	8,12,1,1,13,0,12,13,1,5,22,1,2,22,2,10,23,0,5,23,1,7,23,2,2,
/* out0506_em-eta6-phi25*/	5,12,0,9,12,1,13,12,2,1,21,2,1,22,2,3,
/* out0507_em-eta7-phi25*/	4,11,1,12,11,2,1,12,0,7,21,2,2,
/* out0508_em-eta8-phi25*/	3,11,0,10,11,1,1,11,2,7,
/* out0509_em-eta9-phi25*/	4,3,0,1,10,1,7,10,2,7,11,0,1,
/* out0510_em-eta10-phi25*/	3,2,1,2,10,0,3,10,2,8,
/* out0511_em-eta11-phi25*/	4,2,0,4,2,1,1,9,1,1,9,2,4,
/* out0512_em-eta12-phi25*/	3,1,1,3,2,0,1,9,2,5,
/* out0513_em-eta13-phi25*/	2,1,0,3,1,1,4,
/* out0514_em-eta14-phi25*/	1,1,0,6,
/* out0515_em-eta15-phi25*/	2,0,1,4,1,0,1,
/* out0516_em-eta16-phi25*/	2,0,0,1,0,1,4,
/* out0517_em-eta17-phi25*/	1,0,0,3,
/* out0518_em-eta18-phi25*/	1,0,0,3,
/* out0519_em-eta19-phi25*/	0,
/* out0520_em-eta0-phi26*/	0,
/* out0521_em-eta1-phi26*/	0,
/* out0522_em-eta2-phi26*/	0,
/* out0523_em-eta3-phi26*/	0,
/* out0524_em-eta4-phi26*/	3,6,0,4,13,1,4,13,2,1,
/* out0525_em-eta5-phi26*/	6,5,1,7,6,0,5,6,2,1,13,0,4,13,1,3,13,2,15,
/* out0526_em-eta6-phi26*/	5,4,1,2,5,0,9,5,1,1,12,1,2,12,2,12,
/* out0527_em-eta7-phi26*/	4,4,0,8,4,1,8,11,2,3,12,2,3,
/* out0528_em-eta8-phi26*/	3,3,1,9,4,0,4,11,2,5,
/* out0529_em-eta9-phi26*/	2,3,0,11,3,1,4,
/* out0530_em-eta10-phi26*/	3,2,1,10,3,0,2,10,2,1,
/* out0531_em-eta11-phi26*/	3,2,0,6,2,1,2,2,2,2,
/* out0532_em-eta12-phi26*/	2,1,1,5,2,0,4,
/* out0533_em-eta13-phi26*/	3,1,0,1,1,1,4,1,2,3,
/* out0534_em-eta14-phi26*/	2,1,0,4,1,2,2,
/* out0535_em-eta15-phi26*/	3,0,1,3,0,2,1,1,0,1,
/* out0536_em-eta16-phi26*/	2,0,1,1,0,2,3,
/* out0537_em-eta17-phi26*/	1,0,2,3,
/* out0538_em-eta18-phi26*/	2,0,0,1,0,2,2,
/* out0539_em-eta19-phi26*/	0,
/* out0540_em-eta0-phi27*/	0,
/* out0541_em-eta1-phi27*/	0,
/* out0542_em-eta2-phi27*/	0,
/* out0543_em-eta3-phi27*/	0,
/* out0544_em-eta4-phi27*/	2,6,0,5,6,2,1,
/* out0545_em-eta5-phi27*/	4,5,1,7,5,2,5,6,0,2,6,2,14,
/* out0546_em-eta6-phi27*/	4,4,1,2,5,0,7,5,1,1,5,2,11,
/* out0547_em-eta7-phi27*/	3,4,0,1,4,1,4,4,2,14,
/* out0548_em-eta8-phi27*/	4,3,1,3,3,2,4,4,0,3,4,2,2,
/* out0549_em-eta9-phi27*/	2,3,0,1,3,2,11,
/* out0550_em-eta10-phi27*/	4,2,1,1,2,2,4,3,0,1,3,2,1,
/* out0551_em-eta11-phi27*/	1,2,2,9,
/* out0552_em-eta12-phi27*/	3,1,2,1,2,0,1,2,2,1,
/* out0553_em-eta13-phi27*/	1,1,2,6,
/* out0554_em-eta14-phi27*/	1,1,2,4,
/* out0555_em-eta15-phi27*/	1,0,2,1,
/* out0556_em-eta16-phi27*/	1,0,2,3,
/* out0557_em-eta17-phi27*/	1,0,2,3,
/* out0558_em-eta18-phi27*/	0,
/* out0559_em-eta19-phi27*/	0,
/* out0560_em-eta0-phi28*/	0,
/* out0561_em-eta1-phi28*/	0,
/* out0562_em-eta2-phi28*/	0,
/* out0563_em-eta3-phi28*/	0,
/* out0564_em-eta4-phi28*/	0,
/* out0565_em-eta5-phi28*/	0,
/* out0566_em-eta6-phi28*/	0,
/* out0567_em-eta7-phi28*/	0,
/* out0568_em-eta8-phi28*/	0,
/* out0569_em-eta9-phi28*/	0,
/* out0570_em-eta10-phi28*/	0,
/* out0571_em-eta11-phi28*/	0,
/* out0572_em-eta12-phi28*/	0,
/* out0573_em-eta13-phi28*/	0,
/* out0574_em-eta14-phi28*/	0,
/* out0575_em-eta15-phi28*/	0,
/* out0576_em-eta16-phi28*/	0,
/* out0577_em-eta17-phi28*/	0,
/* out0578_em-eta18-phi28*/	0,
/* out0579_em-eta19-phi28*/	0,
/* out0580_em-eta0-phi29*/	0,
/* out0581_em-eta1-phi29*/	0,
/* out0582_em-eta2-phi29*/	0,
/* out0583_em-eta3-phi29*/	0,
/* out0584_em-eta4-phi29*/	0,
/* out0585_em-eta5-phi29*/	0,
/* out0586_em-eta6-phi29*/	0,
/* out0587_em-eta7-phi29*/	0,
/* out0588_em-eta8-phi29*/	0,
/* out0589_em-eta9-phi29*/	0,
/* out0590_em-eta10-phi29*/	0,
/* out0591_em-eta11-phi29*/	0,
/* out0592_em-eta12-phi29*/	0,
/* out0593_em-eta13-phi29*/	0,
/* out0594_em-eta14-phi29*/	0,
/* out0595_em-eta15-phi29*/	0,
/* out0596_em-eta16-phi29*/	0,
/* out0597_em-eta17-phi29*/	0,
/* out0598_em-eta18-phi29*/	0,
/* out0599_em-eta19-phi29*/	0
};