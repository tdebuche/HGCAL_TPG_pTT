parameter integer matrixH [0:2178] = {
/* num inputs = 133(in0-in132) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 5 */
//* total number of input in adders 849 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	1, 110, 3, 
/* out0002_had-eta2-phi0*/	1, 110, 4, 
/* out0003_had-eta3-phi0*/	2, 109, 3, 110, 1, 
/* out0004_had-eta4-phi0*/	1, 109, 4, 
/* out0005_had-eta5-phi0*/	1, 109, 1, 
/* out0006_had-eta6-phi0*/	1, 63, 1, 
/* out0007_had-eta7-phi0*/	2, 62, 2, 63, 9, 
/* out0008_had-eta8-phi0*/	1, 62, 6, 
/* out0009_had-eta9-phi0*/	2, 61, 3, 62, 1, 
/* out0010_had-eta10-phi0*/	1, 61, 4, 
/* out0011_had-eta11-phi0*/	2, 60, 2, 104, 5, 
/* out0012_had-eta12-phi0*/	2, 60, 3, 104, 5, 
/* out0013_had-eta13-phi0*/	3, 59, 1, 103, 3, 104, 1, 
/* out0014_had-eta14-phi0*/	2, 59, 2, 103, 4, 
/* out0015_had-eta15-phi0*/	3, 59, 1, 102, 1, 103, 2, 
/* out0016_had-eta16-phi0*/	2, 58, 1, 102, 3, 
/* out0017_had-eta17-phi0*/	2, 58, 2, 102, 2, 
/* out0018_had-eta18-phi0*/	1, 102, 2, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	1, 110, 3, 
/* out0022_had-eta2-phi1*/	1, 110, 4, 
/* out0023_had-eta3-phi1*/	2, 109, 3, 110, 1, 
/* out0024_had-eta4-phi1*/	1, 109, 4, 
/* out0025_had-eta5-phi1*/	1, 109, 1, 
/* out0026_had-eta6-phi1*/	2, 57, 1, 63, 1, 
/* out0027_had-eta7-phi1*/	3, 57, 5, 62, 1, 63, 5, 
/* out0028_had-eta8-phi1*/	2, 56, 1, 62, 5, 
/* out0029_had-eta9-phi1*/	3, 56, 1, 61, 4, 62, 1, 
/* out0030_had-eta10-phi1*/	1, 61, 5, 
/* out0031_had-eta11-phi1*/	3, 60, 4, 100, 5, 104, 2, 
/* out0032_had-eta12-phi1*/	3, 60, 4, 98, 2, 104, 3, 
/* out0033_had-eta13-phi1*/	4, 59, 2, 60, 1, 98, 1, 103, 3, 
/* out0034_had-eta14-phi1*/	2, 59, 3, 103, 3, 
/* out0035_had-eta15-phi1*/	4, 59, 2, 97, 1, 102, 1, 103, 1, 
/* out0036_had-eta16-phi1*/	2, 58, 3, 102, 2, 
/* out0037_had-eta17-phi1*/	2, 58, 2, 102, 2, 
/* out0038_had-eta18-phi1*/	1, 102, 1, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	1, 112, 3, 
/* out0042_had-eta2-phi2*/	1, 112, 4, 
/* out0043_had-eta3-phi2*/	2, 111, 3, 112, 1, 
/* out0044_had-eta4-phi2*/	1, 111, 4, 
/* out0045_had-eta5-phi2*/	1, 111, 1, 
/* out0046_had-eta6-phi2*/	1, 57, 1, 
/* out0047_had-eta7-phi2*/	2, 50, 1, 57, 8, 
/* out0048_had-eta8-phi2*/	2, 56, 6, 57, 1, 
/* out0049_had-eta9-phi2*/	2, 55, 1, 56, 5, 
/* out0050_had-eta10-phi2*/	2, 55, 5, 100, 2, 
/* out0051_had-eta11-phi2*/	4, 55, 3, 60, 1, 98, 1, 100, 8, 
/* out0052_had-eta12-phi2*/	3, 54, 2, 60, 1, 98, 4, 
/* out0053_had-eta13-phi2*/	3, 54, 1, 59, 1, 98, 3, 
/* out0054_had-eta14-phi2*/	2, 59, 2, 97, 3, 
/* out0055_had-eta15-phi2*/	2, 59, 2, 97, 2, 
/* out0056_had-eta16-phi2*/	3, 58, 3, 97, 1, 102, 1, 
/* out0057_had-eta17-phi2*/	3, 58, 2, 96, 1, 102, 1, 
/* out0058_had-eta18-phi2*/	1, 96, 1, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 112, 3, 
/* out0062_had-eta2-phi3*/	1, 112, 4, 
/* out0063_had-eta3-phi3*/	2, 111, 3, 112, 1, 
/* out0064_had-eta4-phi3*/	1, 111, 4, 
/* out0065_had-eta5-phi3*/	1, 111, 1, 
/* out0066_had-eta6-phi3*/	1, 52, 1, 
/* out0067_had-eta7-phi3*/	1, 50, 7, 
/* out0068_had-eta8-phi3*/	3, 49, 1, 50, 5, 56, 2, 
/* out0069_had-eta9-phi3*/	3, 49, 4, 55, 1, 56, 1, 
/* out0070_had-eta10-phi3*/	3, 55, 4, 100, 1, 101, 1, 
/* out0071_had-eta11-phi3*/	3, 54, 1, 55, 2, 101, 6, 
/* out0072_had-eta12-phi3*/	4, 54, 4, 98, 3, 99, 1, 101, 1, 
/* out0073_had-eta13-phi3*/	3, 54, 3, 98, 2, 99, 1, 
/* out0074_had-eta14-phi3*/	2, 53, 2, 97, 3, 
/* out0075_had-eta15-phi3*/	2, 53, 2, 97, 3, 
/* out0076_had-eta16-phi3*/	4, 53, 1, 58, 2, 96, 1, 97, 1, 
/* out0077_had-eta17-phi3*/	2, 58, 1, 96, 2, 
/* out0078_had-eta18-phi3*/	1, 96, 2, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 114, 3, 
/* out0082_had-eta2-phi4*/	1, 114, 4, 
/* out0083_had-eta3-phi4*/	2, 113, 3, 114, 1, 
/* out0084_had-eta4-phi4*/	1, 113, 4, 
/* out0085_had-eta5-phi4*/	1, 113, 1, 
/* out0086_had-eta6-phi4*/	1, 52, 5, 
/* out0087_had-eta7-phi4*/	3, 50, 2, 51, 2, 52, 8, 
/* out0088_had-eta8-phi4*/	3, 49, 3, 50, 1, 51, 3, 
/* out0089_had-eta9-phi4*/	1, 49, 6, 
/* out0090_had-eta10-phi4*/	3, 48, 4, 49, 1, 101, 1, 
/* out0091_had-eta11-phi4*/	2, 48, 4, 101, 6, 
/* out0092_had-eta12-phi4*/	4, 48, 1, 54, 3, 99, 3, 101, 1, 
/* out0093_had-eta13-phi4*/	3, 44, 1, 54, 2, 99, 3, 
/* out0094_had-eta14-phi4*/	3, 53, 2, 97, 1, 99, 2, 
/* out0095_had-eta15-phi4*/	3, 53, 2, 92, 1, 97, 1, 
/* out0096_had-eta16-phi4*/	3, 53, 2, 92, 1, 96, 1, 
/* out0097_had-eta17-phi4*/	1, 96, 2, 
/* out0098_had-eta18-phi4*/	1, 96, 2, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 114, 3, 
/* out0102_had-eta2-phi5*/	1, 114, 4, 
/* out0103_had-eta3-phi5*/	2, 113, 3, 114, 1, 
/* out0104_had-eta4-phi5*/	1, 113, 4, 
/* out0105_had-eta5-phi5*/	1, 113, 1, 
/* out0106_had-eta6-phi5*/	2, 52, 1, 70, 2, 
/* out0107_had-eta7-phi5*/	3, 51, 5, 52, 1, 70, 6, 
/* out0108_had-eta8-phi5*/	2, 51, 6, 68, 1, 
/* out0109_had-eta9-phi5*/	2, 49, 1, 68, 5, 
/* out0110_had-eta10-phi5*/	2, 48, 3, 68, 1, 
/* out0111_had-eta11-phi5*/	2, 48, 4, 94, 6, 
/* out0112_had-eta12-phi5*/	3, 44, 3, 94, 2, 99, 2, 
/* out0113_had-eta13-phi5*/	2, 44, 3, 99, 3, 
/* out0114_had-eta14-phi5*/	4, 44, 1, 53, 2, 92, 2, 99, 1, 
/* out0115_had-eta15-phi5*/	2, 53, 2, 92, 2, 
/* out0116_had-eta16-phi5*/	2, 53, 1, 92, 2, 
/* out0117_had-eta17-phi5*/	1, 96, 2, 
/* out0118_had-eta18-phi5*/	1, 96, 2, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 116, 3, 
/* out0122_had-eta2-phi6*/	1, 116, 4, 
/* out0123_had-eta3-phi6*/	2, 115, 3, 116, 1, 
/* out0124_had-eta4-phi6*/	1, 115, 4, 
/* out0125_had-eta5-phi6*/	1, 115, 1, 
/* out0126_had-eta6-phi6*/	2, 70, 2, 71, 1, 
/* out0127_had-eta7-phi6*/	3, 69, 5, 70, 6, 71, 1, 
/* out0128_had-eta8-phi6*/	2, 68, 1, 69, 6, 
/* out0129_had-eta9-phi6*/	2, 46, 1, 68, 6, 
/* out0130_had-eta10-phi6*/	2, 45, 3, 68, 2, 
/* out0131_had-eta11-phi6*/	2, 45, 4, 94, 6, 
/* out0132_had-eta12-phi6*/	3, 44, 3, 93, 2, 94, 2, 
/* out0133_had-eta13-phi6*/	2, 44, 3, 93, 3, 
/* out0134_had-eta14-phi6*/	4, 39, 2, 44, 1, 92, 2, 93, 1, 
/* out0135_had-eta15-phi6*/	2, 39, 2, 92, 2, 
/* out0136_had-eta16-phi6*/	2, 39, 1, 92, 2, 
/* out0137_had-eta17-phi6*/	1, 105, 2, 
/* out0138_had-eta18-phi6*/	1, 105, 2, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 116, 3, 
/* out0142_had-eta2-phi7*/	1, 116, 4, 
/* out0143_had-eta3-phi7*/	2, 115, 3, 116, 1, 
/* out0144_had-eta4-phi7*/	1, 115, 4, 
/* out0145_had-eta5-phi7*/	1, 115, 1, 
/* out0146_had-eta6-phi7*/	1, 71, 5, 
/* out0147_had-eta7-phi7*/	3, 47, 2, 69, 2, 71, 8, 
/* out0148_had-eta8-phi7*/	3, 46, 3, 47, 1, 69, 3, 
/* out0149_had-eta9-phi7*/	1, 46, 6, 
/* out0150_had-eta10-phi7*/	3, 45, 4, 46, 1, 95, 1, 
/* out0151_had-eta11-phi7*/	2, 45, 4, 95, 6, 
/* out0152_had-eta12-phi7*/	4, 40, 3, 45, 1, 93, 3, 95, 1, 
/* out0153_had-eta13-phi7*/	3, 40, 2, 44, 1, 93, 3, 
/* out0154_had-eta14-phi7*/	3, 39, 2, 93, 2, 106, 1, 
/* out0155_had-eta15-phi7*/	3, 39, 2, 92, 1, 106, 1, 
/* out0156_had-eta16-phi7*/	3, 39, 2, 92, 1, 105, 1, 
/* out0157_had-eta17-phi7*/	1, 105, 2, 
/* out0158_had-eta18-phi7*/	1, 105, 2, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 118, 3, 
/* out0162_had-eta2-phi8*/	1, 118, 4, 
/* out0163_had-eta3-phi8*/	2, 117, 3, 118, 1, 
/* out0164_had-eta4-phi8*/	1, 117, 4, 
/* out0165_had-eta5-phi8*/	1, 117, 1, 
/* out0166_had-eta6-phi8*/	1, 71, 1, 
/* out0167_had-eta7-phi8*/	1, 47, 7, 
/* out0168_had-eta8-phi8*/	3, 42, 2, 46, 1, 47, 5, 
/* out0169_had-eta9-phi8*/	3, 41, 1, 42, 1, 46, 4, 
/* out0170_had-eta10-phi8*/	3, 41, 4, 95, 1, 108, 1, 
/* out0171_had-eta11-phi8*/	3, 40, 1, 41, 2, 95, 6, 
/* out0172_had-eta12-phi8*/	4, 40, 4, 93, 1, 95, 1, 107, 3, 
/* out0173_had-eta13-phi8*/	3, 40, 3, 93, 1, 107, 2, 
/* out0174_had-eta14-phi8*/	2, 39, 2, 106, 3, 
/* out0175_had-eta15-phi8*/	2, 39, 2, 106, 3, 
/* out0176_had-eta16-phi8*/	4, 33, 2, 39, 1, 105, 1, 106, 1, 
/* out0177_had-eta17-phi8*/	2, 33, 1, 105, 2, 
/* out0178_had-eta18-phi8*/	1, 105, 2, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 118, 3, 
/* out0182_had-eta2-phi9*/	1, 118, 4, 
/* out0183_had-eta3-phi9*/	2, 117, 3, 118, 1, 
/* out0184_had-eta4-phi9*/	1, 117, 4, 
/* out0185_had-eta5-phi9*/	1, 117, 1, 
/* out0186_had-eta6-phi9*/	1, 43, 1, 
/* out0187_had-eta7-phi9*/	2, 43, 8, 47, 1, 
/* out0188_had-eta8-phi9*/	2, 42, 6, 43, 1, 
/* out0189_had-eta9-phi9*/	2, 41, 1, 42, 5, 
/* out0190_had-eta10-phi9*/	2, 41, 5, 108, 2, 
/* out0191_had-eta11-phi9*/	4, 35, 1, 41, 3, 107, 1, 108, 8, 
/* out0192_had-eta12-phi9*/	3, 35, 1, 40, 2, 107, 4, 
/* out0193_had-eta13-phi9*/	3, 34, 1, 40, 1, 107, 3, 
/* out0194_had-eta14-phi9*/	2, 34, 2, 106, 3, 
/* out0195_had-eta15-phi9*/	2, 34, 2, 106, 2, 
/* out0196_had-eta16-phi9*/	3, 33, 3, 89, 1, 106, 1, 
/* out0197_had-eta17-phi9*/	3, 33, 2, 89, 1, 105, 1, 
/* out0198_had-eta18-phi9*/	1, 105, 1, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 120, 3, 
/* out0202_had-eta2-phi10*/	1, 120, 4, 
/* out0203_had-eta3-phi10*/	2, 119, 3, 120, 1, 
/* out0204_had-eta4-phi10*/	1, 119, 4, 
/* out0205_had-eta5-phi10*/	1, 119, 1, 
/* out0206_had-eta6-phi10*/	2, 38, 1, 43, 1, 
/* out0207_had-eta7-phi10*/	3, 37, 1, 38, 5, 43, 5, 
/* out0208_had-eta8-phi10*/	2, 37, 5, 42, 1, 
/* out0209_had-eta9-phi10*/	3, 36, 4, 37, 1, 42, 1, 
/* out0210_had-eta10-phi10*/	1, 36, 5, 
/* out0211_had-eta11-phi10*/	3, 35, 4, 91, 2, 108, 5, 
/* out0212_had-eta12-phi10*/	3, 35, 4, 91, 2, 107, 2, 
/* out0213_had-eta13-phi10*/	4, 34, 2, 35, 1, 90, 2, 107, 1, 
/* out0214_had-eta14-phi10*/	2, 34, 3, 90, 3, 
/* out0215_had-eta15-phi10*/	4, 34, 2, 89, 1, 90, 1, 106, 1, 
/* out0216_had-eta16-phi10*/	2, 33, 3, 89, 2, 
/* out0217_had-eta17-phi10*/	2, 33, 2, 89, 2, 
/* out0218_had-eta18-phi10*/	1, 89, 1, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 120, 3, 
/* out0222_had-eta2-phi11*/	1, 120, 4, 
/* out0223_had-eta3-phi11*/	2, 119, 3, 120, 1, 
/* out0224_had-eta4-phi11*/	1, 119, 4, 
/* out0225_had-eta5-phi11*/	1, 119, 1, 
/* out0226_had-eta6-phi11*/	1, 38, 1, 
/* out0227_had-eta7-phi11*/	3, 32, 2, 37, 2, 38, 9, 
/* out0228_had-eta8-phi11*/	2, 32, 1, 37, 6, 
/* out0229_had-eta9-phi11*/	3, 31, 2, 36, 3, 37, 1, 
/* out0230_had-eta10-phi11*/	2, 30, 1, 36, 4, 
/* out0231_had-eta11-phi11*/	3, 30, 2, 35, 2, 91, 4, 
/* out0232_had-eta12-phi11*/	3, 29, 1, 35, 3, 91, 4, 
/* out0233_had-eta13-phi11*/	4, 29, 1, 34, 1, 90, 3, 91, 1, 
/* out0234_had-eta14-phi11*/	2, 34, 2, 90, 3, 
/* out0235_had-eta15-phi11*/	4, 28, 1, 34, 1, 89, 1, 90, 2, 
/* out0236_had-eta16-phi11*/	3, 28, 1, 33, 1, 89, 2, 
/* out0237_had-eta17-phi11*/	2, 33, 2, 89, 2, 
/* out0238_had-eta18-phi11*/	1, 89, 1, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 122, 3, 
/* out0242_had-eta2-phi12*/	1, 122, 4, 
/* out0243_had-eta3-phi12*/	2, 121, 3, 122, 1, 
/* out0244_had-eta4-phi12*/	1, 121, 4, 
/* out0245_had-eta5-phi12*/	1, 121, 1, 
/* out0246_had-eta6-phi12*/	0, 
/* out0247_had-eta7-phi12*/	1, 32, 9, 
/* out0248_had-eta8-phi12*/	2, 31, 4, 32, 3, 
/* out0249_had-eta9-phi12*/	1, 31, 6, 
/* out0250_had-eta10-phi12*/	2, 30, 4, 31, 1, 
/* out0251_had-eta11-phi12*/	3, 30, 4, 88, 6, 91, 1, 
/* out0252_had-eta12-phi12*/	4, 29, 3, 30, 1, 87, 2, 91, 2, 
/* out0253_had-eta13-phi12*/	3, 29, 3, 87, 3, 90, 1, 
/* out0254_had-eta14-phi12*/	4, 28, 1, 29, 2, 86, 1, 90, 1, 
/* out0255_had-eta15-phi12*/	2, 28, 2, 86, 2, 
/* out0256_had-eta16-phi12*/	3, 28, 2, 86, 1, 89, 1, 
/* out0257_had-eta17-phi12*/	3, 28, 1, 85, 1, 89, 1, 
/* out0258_had-eta18-phi12*/	1, 85, 2, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 122, 3, 
/* out0262_had-eta2-phi13*/	1, 122, 4, 
/* out0263_had-eta3-phi13*/	2, 121, 3, 122, 1, 
/* out0264_had-eta4-phi13*/	1, 121, 4, 
/* out0265_had-eta5-phi13*/	1, 121, 1, 
/* out0266_had-eta6-phi13*/	1, 27, 2, 
/* out0267_had-eta7-phi13*/	3, 26, 3, 27, 9, 32, 1, 
/* out0268_had-eta8-phi13*/	2, 26, 6, 31, 1, 
/* out0269_had-eta9-phi13*/	2, 25, 3, 31, 2, 
/* out0270_had-eta10-phi13*/	2, 25, 3, 30, 2, 
/* out0271_had-eta11-phi13*/	3, 24, 2, 30, 2, 88, 9, 
/* out0272_had-eta12-phi13*/	3, 24, 1, 29, 2, 87, 4, 
/* out0273_had-eta13-phi13*/	2, 29, 3, 87, 4, 
/* out0274_had-eta14-phi13*/	5, 23, 1, 28, 1, 29, 1, 86, 2, 87, 1, 
/* out0275_had-eta15-phi13*/	2, 28, 2, 86, 3, 
/* out0276_had-eta16-phi13*/	2, 28, 2, 86, 2, 
/* out0277_had-eta17-phi13*/	2, 28, 1, 85, 3, 
/* out0278_had-eta18-phi13*/	1, 85, 2, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 124, 3, 
/* out0282_had-eta2-phi14*/	1, 124, 4, 
/* out0283_had-eta3-phi14*/	2, 123, 3, 124, 1, 
/* out0284_had-eta4-phi14*/	1, 123, 4, 
/* out0285_had-eta5-phi14*/	1, 123, 1, 
/* out0286_had-eta6-phi14*/	2, 21, 2, 27, 2, 
/* out0287_had-eta7-phi14*/	3, 21, 7, 26, 2, 27, 3, 
/* out0288_had-eta8-phi14*/	2, 19, 2, 26, 5, 
/* out0289_had-eta9-phi14*/	2, 19, 1, 25, 5, 
/* out0290_had-eta10-phi14*/	3, 24, 1, 25, 4, 84, 1, 
/* out0291_had-eta11-phi14*/	3, 24, 4, 84, 5, 88, 1, 
/* out0292_had-eta12-phi14*/	3, 24, 3, 84, 3, 87, 1, 
/* out0293_had-eta13-phi14*/	3, 23, 3, 82, 2, 87, 1, 
/* out0294_had-eta14-phi14*/	3, 23, 2, 82, 1, 86, 1, 
/* out0295_had-eta15-phi14*/	3, 23, 1, 28, 1, 86, 2, 
/* out0296_had-eta16-phi14*/	3, 22, 1, 28, 1, 86, 2, 
/* out0297_had-eta17-phi14*/	2, 22, 1, 85, 3, 
/* out0298_had-eta18-phi14*/	1, 85, 2, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 124, 3, 
/* out0302_had-eta2-phi15*/	1, 124, 4, 
/* out0303_had-eta3-phi15*/	2, 123, 3, 124, 1, 
/* out0304_had-eta4-phi15*/	1, 123, 4, 
/* out0305_had-eta5-phi15*/	1, 123, 1, 
/* out0306_had-eta6-phi15*/	0, 
/* out0307_had-eta7-phi15*/	2, 20, 2, 21, 7, 
/* out0308_had-eta8-phi15*/	1, 19, 7, 
/* out0309_had-eta9-phi15*/	3, 17, 2, 19, 4, 25, 1, 
/* out0310_had-eta10-phi15*/	2, 17, 5, 84, 1, 
/* out0311_had-eta11-phi15*/	4, 16, 1, 17, 1, 24, 3, 84, 4, 
/* out0312_had-eta12-phi15*/	4, 16, 1, 24, 2, 82, 1, 84, 2, 
/* out0313_had-eta13-phi15*/	2, 23, 3, 82, 4, 
/* out0314_had-eta14-phi15*/	2, 23, 3, 82, 3, 
/* out0315_had-eta15-phi15*/	3, 22, 1, 23, 1, 81, 2, 
/* out0316_had-eta16-phi15*/	2, 22, 2, 81, 2, 
/* out0317_had-eta17-phi15*/	3, 22, 2, 81, 1, 85, 2, 
/* out0318_had-eta18-phi15*/	1, 85, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 126, 3, 
/* out0322_had-eta2-phi16*/	1, 126, 4, 
/* out0323_had-eta3-phi16*/	2, 125, 3, 126, 1, 
/* out0324_had-eta4-phi16*/	1, 125, 4, 
/* out0325_had-eta5-phi16*/	1, 125, 1, 
/* out0326_had-eta6-phi16*/	1, 20, 1, 
/* out0327_had-eta7-phi16*/	1, 20, 9, 
/* out0328_had-eta8-phi16*/	3, 18, 3, 19, 1, 20, 2, 
/* out0329_had-eta9-phi16*/	3, 17, 2, 18, 3, 19, 1, 
/* out0330_had-eta10-phi16*/	1, 17, 5, 
/* out0331_had-eta11-phi16*/	3, 16, 3, 17, 1, 83, 4, 
/* out0332_had-eta12-phi16*/	2, 16, 3, 83, 4, 
/* out0333_had-eta13-phi16*/	4, 16, 2, 23, 1, 82, 3, 83, 1, 
/* out0334_had-eta14-phi16*/	4, 11, 1, 23, 1, 79, 1, 82, 2, 
/* out0335_had-eta15-phi16*/	3, 11, 1, 22, 1, 81, 2, 
/* out0336_had-eta16-phi16*/	2, 22, 2, 81, 2, 
/* out0337_had-eta17-phi16*/	2, 22, 2, 81, 2, 
/* out0338_had-eta18-phi16*/	0, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 126, 3, 
/* out0342_had-eta2-phi17*/	1, 126, 4, 
/* out0343_had-eta3-phi17*/	2, 125, 3, 126, 1, 
/* out0344_had-eta4-phi17*/	1, 125, 4, 
/* out0345_had-eta5-phi17*/	1, 125, 1, 
/* out0346_had-eta6-phi17*/	0, 
/* out0347_had-eta7-phi17*/	2, 20, 2, 67, 6, 
/* out0348_had-eta8-phi17*/	2, 18, 5, 67, 2, 
/* out0349_had-eta9-phi17*/	2, 18, 5, 64, 1, 
/* out0350_had-eta10-phi17*/	1, 64, 5, 
/* out0351_had-eta11-phi17*/	3, 16, 2, 64, 2, 83, 3, 
/* out0352_had-eta12-phi17*/	2, 16, 3, 83, 4, 
/* out0353_had-eta13-phi17*/	3, 11, 2, 16, 1, 79, 3, 
/* out0354_had-eta14-phi17*/	2, 11, 2, 79, 3, 
/* out0355_had-eta15-phi17*/	3, 11, 2, 79, 1, 81, 2, 
/* out0356_had-eta16-phi17*/	2, 22, 2, 81, 2, 
/* out0357_had-eta17-phi17*/	2, 22, 2, 81, 1, 
/* out0358_had-eta18-phi17*/	0, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 128, 3, 
/* out0362_had-eta2-phi18*/	1, 128, 4, 
/* out0363_had-eta3-phi18*/	2, 127, 3, 128, 1, 
/* out0364_had-eta4-phi18*/	1, 127, 4, 
/* out0365_had-eta5-phi18*/	1, 127, 1, 
/* out0366_had-eta6-phi18*/	0, 
/* out0367_had-eta7-phi18*/	2, 66, 2, 67, 6, 
/* out0368_had-eta8-phi18*/	2, 65, 5, 67, 2, 
/* out0369_had-eta9-phi18*/	2, 64, 1, 65, 5, 
/* out0370_had-eta10-phi18*/	1, 64, 5, 
/* out0371_had-eta11-phi18*/	3, 12, 2, 64, 2, 80, 3, 
/* out0372_had-eta12-phi18*/	2, 12, 3, 80, 4, 
/* out0373_had-eta13-phi18*/	3, 11, 2, 12, 1, 79, 3, 
/* out0374_had-eta14-phi18*/	2, 11, 2, 79, 3, 
/* out0375_had-eta15-phi18*/	3, 11, 2, 76, 2, 79, 1, 
/* out0376_had-eta16-phi18*/	2, 5, 2, 76, 2, 
/* out0377_had-eta17-phi18*/	2, 5, 2, 76, 1, 
/* out0378_had-eta18-phi18*/	0, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 128, 3, 
/* out0382_had-eta2-phi19*/	1, 128, 4, 
/* out0383_had-eta3-phi19*/	2, 127, 3, 128, 1, 
/* out0384_had-eta4-phi19*/	1, 127, 4, 
/* out0385_had-eta5-phi19*/	1, 127, 1, 
/* out0386_had-eta6-phi19*/	1, 66, 1, 
/* out0387_had-eta7-phi19*/	1, 66, 9, 
/* out0388_had-eta8-phi19*/	3, 14, 1, 65, 3, 66, 2, 
/* out0389_had-eta9-phi19*/	3, 13, 2, 14, 1, 65, 3, 
/* out0390_had-eta10-phi19*/	1, 13, 5, 
/* out0391_had-eta11-phi19*/	3, 12, 3, 13, 1, 80, 4, 
/* out0392_had-eta12-phi19*/	2, 12, 3, 80, 4, 
/* out0393_had-eta13-phi19*/	4, 6, 1, 12, 2, 77, 3, 80, 1, 
/* out0394_had-eta14-phi19*/	4, 6, 1, 11, 1, 77, 2, 79, 1, 
/* out0395_had-eta15-phi19*/	3, 5, 1, 11, 1, 76, 2, 
/* out0396_had-eta16-phi19*/	2, 5, 2, 76, 2, 
/* out0397_had-eta17-phi19*/	2, 5, 2, 76, 2, 
/* out0398_had-eta18-phi19*/	0, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 130, 3, 
/* out0402_had-eta2-phi20*/	1, 130, 4, 
/* out0403_had-eta3-phi20*/	2, 129, 3, 130, 1, 
/* out0404_had-eta4-phi20*/	1, 129, 4, 
/* out0405_had-eta5-phi20*/	1, 129, 1, 
/* out0406_had-eta6-phi20*/	0, 
/* out0407_had-eta7-phi20*/	2, 15, 7, 66, 2, 
/* out0408_had-eta8-phi20*/	1, 14, 7, 
/* out0409_had-eta9-phi20*/	3, 8, 1, 13, 2, 14, 4, 
/* out0410_had-eta10-phi20*/	2, 13, 5, 78, 1, 
/* out0411_had-eta11-phi20*/	4, 7, 3, 12, 1, 13, 1, 78, 4, 
/* out0412_had-eta12-phi20*/	4, 7, 2, 12, 1, 77, 1, 78, 2, 
/* out0413_had-eta13-phi20*/	2, 6, 3, 77, 4, 
/* out0414_had-eta14-phi20*/	2, 6, 3, 77, 3, 
/* out0415_had-eta15-phi20*/	3, 5, 1, 6, 1, 76, 2, 
/* out0416_had-eta16-phi20*/	2, 5, 2, 76, 2, 
/* out0417_had-eta17-phi20*/	3, 5, 2, 72, 2, 76, 1, 
/* out0418_had-eta18-phi20*/	1, 72, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 130, 3, 
/* out0422_had-eta2-phi21*/	1, 130, 4, 
/* out0423_had-eta3-phi21*/	2, 129, 3, 130, 1, 
/* out0424_had-eta4-phi21*/	1, 129, 4, 
/* out0425_had-eta5-phi21*/	1, 129, 1, 
/* out0426_had-eta6-phi21*/	2, 10, 2, 15, 2, 
/* out0427_had-eta7-phi21*/	3, 9, 2, 10, 3, 15, 7, 
/* out0428_had-eta8-phi21*/	2, 9, 5, 14, 2, 
/* out0429_had-eta9-phi21*/	2, 8, 5, 14, 1, 
/* out0430_had-eta10-phi21*/	3, 7, 1, 8, 4, 78, 1, 
/* out0431_had-eta11-phi21*/	3, 7, 4, 75, 1, 78, 5, 
/* out0432_had-eta12-phi21*/	3, 7, 3, 74, 1, 78, 3, 
/* out0433_had-eta13-phi21*/	3, 6, 3, 74, 1, 77, 2, 
/* out0434_had-eta14-phi21*/	3, 6, 2, 73, 1, 77, 1, 
/* out0435_had-eta15-phi21*/	3, 0, 1, 6, 1, 73, 2, 
/* out0436_had-eta16-phi21*/	3, 0, 1, 5, 1, 73, 2, 
/* out0437_had-eta17-phi21*/	2, 5, 1, 72, 3, 
/* out0438_had-eta18-phi21*/	1, 72, 2, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 132, 3, 
/* out0442_had-eta2-phi22*/	1, 132, 4, 
/* out0443_had-eta3-phi22*/	2, 131, 3, 132, 1, 
/* out0444_had-eta4-phi22*/	1, 131, 4, 
/* out0445_had-eta5-phi22*/	1, 131, 1, 
/* out0446_had-eta6-phi22*/	1, 10, 2, 
/* out0447_had-eta7-phi22*/	3, 4, 2, 9, 3, 10, 9, 
/* out0448_had-eta8-phi22*/	2, 3, 1, 9, 6, 
/* out0449_had-eta9-phi22*/	2, 3, 2, 8, 3, 
/* out0450_had-eta10-phi22*/	2, 2, 2, 8, 3, 
/* out0451_had-eta11-phi22*/	3, 2, 3, 7, 2, 75, 9, 
/* out0452_had-eta12-phi22*/	3, 1, 3, 7, 1, 74, 4, 
/* out0453_had-eta13-phi22*/	2, 1, 3, 74, 4, 
/* out0454_had-eta14-phi22*/	5, 0, 1, 1, 1, 6, 1, 73, 2, 74, 1, 
/* out0455_had-eta15-phi22*/	2, 0, 3, 73, 3, 
/* out0456_had-eta16-phi22*/	2, 0, 2, 73, 2, 
/* out0457_had-eta17-phi22*/	2, 0, 1, 72, 3, 
/* out0458_had-eta18-phi22*/	1, 72, 2, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 132, 3, 
/* out0462_had-eta2-phi23*/	1, 132, 4, 
/* out0463_had-eta3-phi23*/	2, 131, 3, 132, 1, 
/* out0464_had-eta4-phi23*/	1, 131, 4, 
/* out0465_had-eta5-phi23*/	1, 131, 1, 
/* out0466_had-eta6-phi23*/	0, 
/* out0467_had-eta7-phi23*/	1, 4, 10, 
/* out0468_had-eta8-phi23*/	2, 3, 5, 4, 4, 
/* out0469_had-eta9-phi23*/	1, 3, 7, 
/* out0470_had-eta10-phi23*/	2, 2, 5, 3, 1, 
/* out0471_had-eta11-phi23*/	2, 2, 5, 75, 6, 
/* out0472_had-eta12-phi23*/	3, 1, 3, 2, 1, 74, 2, 
/* out0473_had-eta13-phi23*/	2, 1, 4, 74, 3, 
/* out0474_had-eta14-phi23*/	3, 0, 1, 1, 2, 73, 1, 
/* out0475_had-eta15-phi23*/	2, 0, 2, 73, 2, 
/* out0476_had-eta16-phi23*/	2, 0, 2, 73, 1, 
/* out0477_had-eta17-phi23*/	2, 0, 2, 72, 1, 
/* out0478_had-eta18-phi23*/	1, 72, 2, 
/* out0479_had-eta19-phi23*/	0, 
};