parameter integer matrixH [0:6827] = {
/* num inputs = 140(in0-in139) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2115 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	4,60,0,1,60,1,3,77,0,10,77,1,15,
/* out0004_em-eta4-phi0*/	2,59,1,7,60,0,7,
/* out0005_em-eta5-phi0*/	3,59,0,15,59,1,6,59,2,5,
/* out0006_em-eta6-phi0*/	3,40,0,3,59,0,1,59,2,1,
/* out0007_em-eta7-phi0*/	2,39,0,2,39,1,10,
/* out0008_em-eta8-phi0*/	1,39,0,13,
/* out0009_em-eta9-phi0*/	1,39,0,1,
/* out0010_em-eta10-phi0*/	2,19,0,1,19,1,5,
/* out0011_em-eta11-phi0*/	5,19,0,15,19,1,5,19,2,7,19,3,7,131,2,10,
/* out0012_em-eta12-phi0*/	8,19,2,2,19,3,9,20,3,13,20,4,2,124,0,3,124,1,2,131,1,2,131,2,2,
/* out0013_em-eta13-phi0*/	2,20,2,1,124,0,9,
/* out0014_em-eta14-phi0*/	3,117,0,1,124,0,2,124,2,1,
/* out0015_em-eta15-phi0*/	1,117,0,5,
/* out0016_em-eta16-phi0*/	3,0,1,4,1,1,8,117,0,4,
/* out0017_em-eta17-phi0*/	4,0,0,1,0,1,11,111,2,1,117,0,1,
/* out0018_em-eta18-phi0*/	2,0,0,10,111,2,3,
/* out0019_em-eta19-phi0*/	2,0,0,2,111,0,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	3,61,1,1,61,2,10,77,0,1,
/* out0023_em-eta3-phi1*/	8,42,0,1,60,1,11,60,2,2,61,0,5,61,1,15,61,2,4,77,0,5,77,1,1,
/* out0024_em-eta4-phi1*/	5,41,0,6,59,1,2,60,0,8,60,1,2,60,2,14,
/* out0025_em-eta5-phi1*/	6,40,0,2,40,1,2,41,0,8,41,2,3,59,1,1,59,2,10,
/* out0026_em-eta6-phi1*/	3,40,0,11,40,1,6,40,2,6,
/* out0027_em-eta7-phi1*/	4,22,0,2,39,1,6,39,2,4,40,2,7,
/* out0028_em-eta8-phi1*/	3,21,1,2,22,0,1,39,2,12,
/* out0029_em-eta9-phi1*/	2,21,0,7,21,1,5,
/* out0030_em-eta10-phi1*/	4,19,1,4,19,4,2,20,1,11,21,0,5,
/* out0031_em-eta11-phi1*/	9,19,1,2,19,2,7,19,4,2,19,5,1,20,0,16,20,1,5,20,4,2,131,1,9,131,2,4,
/* out0032_em-eta12-phi1*/	7,20,2,8,20,3,3,20,4,12,20,5,6,124,1,9,131,1,4,132,0,1,
/* out0033_em-eta13-phi1*/	5,2,0,9,20,2,7,124,0,2,124,1,3,124,2,5,
/* out0034_em-eta14-phi1*/	4,2,0,1,2,3,5,117,1,4,124,2,5,
/* out0035_em-eta15-phi1*/	4,0,4,8,2,3,1,117,0,3,117,1,5,
/* out0036_em-eta16-phi1*/	5,0,4,2,1,0,4,1,1,8,117,0,2,117,2,4,
/* out0037_em-eta17-phi1*/	5,0,1,1,0,2,8,1,0,3,111,2,4,117,2,2,
/* out0038_em-eta18-phi1*/	5,0,0,2,0,2,4,0,3,4,111,0,2,111,2,4,
/* out0039_em-eta19-phi1*/	3,0,0,1,0,3,5,111,0,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	3,43,1,7,61,0,3,61,2,2,
/* out0043_em-eta3-phi2*/	5,42,0,10,42,1,11,43,0,7,43,1,6,61,0,8,
/* out0044_em-eta4-phi2*/	6,24,0,1,24,1,1,41,0,1,41,1,10,42,0,5,42,2,14,
/* out0045_em-eta5-phi2*/	6,23,1,5,24,0,1,40,1,1,41,0,1,41,1,6,41,2,13,
/* out0046_em-eta6-phi2*/	5,22,1,1,23,0,10,23,1,1,40,1,7,40,2,2,
/* out0047_em-eta7-phi2*/	4,22,0,11,22,1,5,22,2,1,40,2,1,
/* out0048_em-eta8-phi2*/	3,21,1,4,22,0,2,22,2,8,
/* out0049_em-eta9-phi2*/	3,21,0,1,21,1,5,21,2,7,
/* out0050_em-eta10-phi2*/	5,4,1,1,5,1,7,19,4,3,21,0,3,21,2,5,
/* out0051_em-eta11-phi2*/	7,4,0,4,4,1,10,19,4,9,19,5,11,131,1,1,132,0,6,132,1,7,
/* out0052_em-eta12-phi2*/	8,2,1,8,3,1,2,4,0,3,19,5,4,20,5,10,124,1,1,132,0,9,132,2,2,
/* out0053_em-eta13-phi2*/	9,2,0,6,2,1,8,2,2,9,2,3,1,124,1,1,124,2,4,125,0,4,125,1,1,132,2,1,
/* out0054_em-eta14-phi2*/	7,2,2,5,2,3,9,3,3,5,3,4,3,117,1,2,124,2,1,125,0,6,
/* out0055_em-eta15-phi2*/	5,0,4,5,0,5,3,3,3,8,117,1,5,117,2,2,
/* out0056_em-eta16-phi2*/	5,0,4,1,0,5,6,1,0,6,1,4,1,117,2,6,
/* out0057_em-eta17-phi2*/	6,0,2,2,1,0,3,1,4,8,111,0,2,111,2,3,117,2,1,
/* out0058_em-eta18-phi2*/	6,0,2,2,0,3,2,1,3,3,1,4,3,111,0,5,111,2,1,
/* out0059_em-eta19-phi2*/	2,0,3,5,1,3,3,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	1,43,1,1,
/* out0063_em-eta3-phi3*/	6,25,0,11,25,1,14,25,2,2,42,1,4,43,0,9,43,1,2,
/* out0064_em-eta4-phi3*/	6,24,0,4,24,1,15,24,2,5,25,0,5,42,1,1,42,2,2,
/* out0065_em-eta5-phi3*/	5,8,0,1,23,1,8,23,2,2,24,0,10,24,2,4,
/* out0066_em-eta6-phi3*/	4,7,1,2,23,0,6,23,1,2,23,2,13,
/* out0067_em-eta7-phi3*/	4,7,0,5,7,1,1,22,1,10,22,2,1,
/* out0068_em-eta8-phi3*/	3,6,0,8,6,1,1,22,2,6,
/* out0069_em-eta9-phi3*/	3,6,0,7,6,2,3,21,2,3,
/* out0070_em-eta10-phi3*/	5,4,4,16,4,5,4,5,0,9,5,1,8,21,2,1,
/* out0071_em-eta11-phi3*/	12,4,0,3,4,1,5,4,2,16,4,3,3,5,0,5,5,1,1,5,4,2,132,1,9,132,2,2,137,0,10,137,1,7,137,2,3,
/* out0072_em-eta12-phi3*/	7,2,4,4,3,1,10,4,0,6,4,3,9,125,1,1,132,2,11,133,0,1,
/* out0073_em-eta13-phi3*/	7,2,2,2,2,4,2,2,5,1,3,0,15,3,1,4,125,0,1,125,1,10,
/* out0074_em-eta14-phi3*/	7,3,0,1,3,2,1,3,3,2,3,4,13,3,5,3,125,0,4,125,2,4,
/* out0075_em-eta15-phi3*/	9,0,5,3,3,2,12,3,3,1,26,1,1,117,2,1,118,0,1,118,1,3,125,0,1,125,2,2,
/* out0076_em-eta16-phi3*/	4,0,5,4,1,4,1,1,5,10,118,0,6,
/* out0077_em-eta17-phi3*/	5,1,2,4,1,4,3,1,5,5,111,0,1,118,0,4,
/* out0078_em-eta18-phi3*/	3,1,2,4,1,3,6,111,0,4,
/* out0079_em-eta19-phi3*/	5,1,3,4,11,1,1,11,5,2,12,1,2,12,5,4,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	1,10,2,5,
/* out0083_em-eta3-phi4*/	5,9,1,5,10,1,14,10,2,10,25,1,2,25,2,12,
/* out0084_em-eta4-phi4*/	5,9,0,15,9,1,9,9,2,1,24,2,5,25,2,2,
/* out0085_em-eta5-phi4*/	4,8,0,6,8,1,15,8,2,3,24,2,2,
/* out0086_em-eta6-phi4*/	5,7,1,10,7,2,1,8,0,9,8,2,1,23,2,1,
/* out0087_em-eta7-phi4*/	3,7,0,9,7,1,3,7,2,7,
/* out0088_em-eta8-phi4*/	3,6,0,1,6,1,12,7,0,2,
/* out0089_em-eta9-phi4*/	2,6,1,1,6,2,10,
/* out0090_em-eta10-phi4*/	7,4,5,12,5,0,2,5,2,1,5,4,2,5,5,13,6,2,1,62,0,2,
/* out0091_em-eta11-phi4*/	9,5,2,11,5,3,8,5,4,12,5,5,3,133,0,1,133,1,6,137,0,6,137,1,9,137,2,13,
/* out0092_em-eta12-phi4*/	8,2,4,4,4,3,4,5,3,8,44,0,12,44,1,1,133,0,11,133,1,2,133,2,1,
/* out0093_em-eta13-phi4*/	9,2,4,6,2,5,11,44,0,3,44,3,4,125,1,4,125,2,2,126,0,1,133,0,3,133,2,1,
/* out0094_em-eta14-phi4*/	5,2,5,4,3,5,13,26,4,3,125,2,7,126,0,2,
/* out0095_em-eta15-phi4*/	6,3,2,3,26,1,1,26,4,1,27,1,13,118,1,6,125,2,1,
/* out0096_em-eta16-phi4*/	6,1,5,1,26,0,1,26,1,12,118,0,2,118,1,3,118,2,2,
/* out0097_em-eta17-phi4*/	4,1,2,5,26,0,6,118,0,2,118,2,3,
/* out0098_em-eta18-phi4*/	5,1,2,3,12,2,8,12,5,2,118,0,1,118,2,1,
/* out0099_em-eta19-phi4*/	5,11,1,5,11,5,10,12,1,10,12,4,1,12,5,9,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	5,9,1,1,9,2,1,10,1,2,10,2,1,114,1,1,
/* out0104_em-eta4-phi5*/	6,9,0,1,9,1,1,9,2,14,102,1,10,114,1,2,114,2,3,
/* out0105_em-eta5-phi5*/	6,8,1,1,8,2,9,90,0,1,90,1,2,102,0,12,102,1,2,
/* out0106_em-eta6-phi5*/	5,7,2,2,8,2,3,90,0,14,90,1,2,90,2,1,
/* out0107_em-eta7-phi5*/	5,7,2,6,78,0,5,78,1,4,90,0,1,90,2,3,
/* out0108_em-eta8-phi5*/	3,6,1,1,78,0,11,78,2,3,
/* out0109_em-eta9-phi5*/	5,6,1,1,6,2,2,62,0,5,62,1,4,78,2,1,
/* out0110_em-eta10-phi5*/	2,62,0,8,62,2,2,
/* out0111_em-eta11-phi5*/	9,5,2,4,44,1,6,45,1,11,62,0,1,62,2,2,133,1,6,138,0,12,138,1,8,138,2,4,
/* out0112_em-eta12-phi5*/	8,44,0,1,44,1,9,44,2,12,44,3,1,45,0,4,45,1,1,133,1,2,133,2,11,
/* out0113_em-eta13-phi5*/	7,44,2,4,44,3,10,45,3,7,45,4,4,126,0,1,126,1,7,133,2,3,
/* out0114_em-eta14-phi5*/	6,26,4,11,26,5,3,44,3,1,45,3,5,126,0,8,126,1,1,
/* out0115_em-eta15-phi5*/	6,26,4,1,26,5,1,27,0,12,27,1,3,118,1,3,126,0,4,
/* out0116_em-eta16-phi5*/	4,26,1,2,26,2,12,118,1,1,118,2,5,
/* out0117_em-eta17-phi5*/	3,26,0,8,26,3,4,118,2,5,
/* out0118_em-eta18-phi5*/	5,12,2,8,12,3,4,12,4,2,12,5,1,26,0,1,
/* out0119_em-eta19-phi5*/	5,11,1,8,11,2,4,11,5,4,12,1,4,12,4,9,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	5,114,1,13,114,2,3,115,1,2,125,1,2,125,2,12,
/* out0124_em-eta4-phi6*/	5,102,1,4,102,2,6,114,2,10,115,0,8,115,1,7,
/* out0125_em-eta5-phi6*/	5,90,1,3,102,0,4,102,2,10,103,0,3,103,1,7,
/* out0126_em-eta6-phi6*/	4,90,1,9,90,2,8,91,1,2,103,0,3,
/* out0127_em-eta7-phi6*/	4,78,1,8,90,2,4,91,0,3,91,1,3,
/* out0128_em-eta8-phi6*/	3,78,1,4,78,2,10,79,0,1,
/* out0129_em-eta9-phi6*/	3,62,1,8,78,2,2,79,0,2,
/* out0130_em-eta10-phi6*/	2,62,1,3,62,2,8,
/* out0131_em-eta11-phi6*/	8,44,4,14,45,1,3,62,2,3,63,0,4,134,1,6,138,0,4,138,1,8,138,2,12,
/* out0132_em-eta12-phi6*/	8,44,4,2,44,5,8,45,0,12,45,1,1,45,4,5,45,5,2,134,0,11,134,1,2,
/* out0133_em-eta13-phi6*/	7,45,2,8,45,3,3,45,4,7,45,5,5,126,1,7,126,2,1,134,0,3,
/* out0134_em-eta14-phi6*/	6,26,5,11,27,5,4,45,2,5,45,3,1,126,1,1,126,2,8,
/* out0135_em-eta15-phi6*/	6,26,5,1,27,0,4,27,4,8,27,5,4,119,1,3,126,2,4,
/* out0136_em-eta16-phi6*/	5,26,2,4,27,3,2,27,4,8,119,0,5,119,1,1,
/* out0137_em-eta17-phi6*/	3,26,3,10,27,3,2,119,0,5,
/* out0138_em-eta18-phi6*/	5,11,2,2,11,3,3,12,3,11,12,4,3,26,3,1,
/* out0139_em-eta19-phi6*/	5,11,0,5,11,1,2,11,2,10,11,3,2,12,4,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	6,115,1,3,115,2,1,125,1,14,125,2,4,126,0,12,126,1,2,
/* out0144_em-eta4-phi7*/	5,115,0,8,115,1,4,115,2,15,116,0,5,126,0,2,
/* out0145_em-eta5-phi7*/	4,103,0,3,103,1,9,103,2,12,116,0,2,
/* out0146_em-eta6-phi7*/	4,91,1,8,91,2,3,103,0,7,103,2,2,
/* out0147_em-eta7-phi7*/	3,91,0,10,91,1,3,91,2,5,
/* out0148_em-eta8-phi7*/	3,79,0,5,79,1,8,91,0,3,
/* out0149_em-eta9-phi7*/	2,79,0,8,79,2,5,
/* out0150_em-eta10-phi7*/	8,62,1,1,62,2,1,63,0,1,63,1,13,63,2,2,64,0,2,64,1,12,79,2,1,
/* out0151_em-eta11-phi7*/	9,63,0,11,63,1,3,63,2,12,63,3,8,134,1,6,134,2,1,139,0,13,139,1,9,139,2,6,
/* out0152_em-eta12-phi7*/	9,44,5,8,45,5,4,46,1,2,47,1,2,63,3,8,64,3,4,134,0,1,134,1,2,134,2,11,
/* out0153_em-eta13-phi7*/	9,45,2,3,45,5,5,46,0,5,46,1,12,126,2,1,127,0,2,127,1,4,134,0,1,134,2,3,
/* out0154_em-eta14-phi7*/	6,27,5,3,46,0,11,46,2,1,46,3,5,126,2,2,127,0,7,
/* out0155_em-eta15-phi7*/	5,27,2,9,27,5,5,46,3,3,119,1,6,127,0,1,
/* out0156_em-eta16-phi7*/	6,27,2,6,27,3,6,28,1,1,119,0,2,119,1,3,119,2,2,
/* out0157_em-eta17-phi7*/	5,26,3,1,27,3,6,28,0,5,119,0,3,119,2,2,
/* out0158_em-eta18-phi7*/	5,11,3,10,12,3,1,28,0,3,119,0,1,119,2,1,
/* out0159_em-eta19-phi7*/	2,11,0,8,11,3,1,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	1,134,2,1,
/* out0163_em-eta3-phi8*/	6,126,0,2,126,1,14,126,2,11,127,0,4,134,0,9,134,2,2,
/* out0164_em-eta4-phi8*/	5,116,0,5,116,1,15,116,2,4,126,2,5,127,0,3,
/* out0165_em-eta5-phi8*/	5,103,2,2,104,1,10,104,2,1,116,0,4,116,2,10,
/* out0166_em-eta6-phi8*/	4,91,2,2,104,0,13,104,1,6,104,2,1,
/* out0167_em-eta7-phi8*/	3,91,2,6,92,0,1,92,1,10,
/* out0168_em-eta8-phi8*/	3,79,1,8,79,2,1,92,0,6,
/* out0169_em-eta9-phi8*/	2,79,2,9,80,1,3,
/* out0170_em-eta10-phi8*/	5,63,4,16,63,5,8,64,0,9,64,1,4,80,0,1,
/* out0171_em-eta11-phi8*/	12,63,2,2,63,5,1,64,0,5,64,2,3,64,3,3,64,4,16,64,5,5,135,0,2,135,1,9,139,0,3,139,1,7,139,2,10,
/* out0172_em-eta12-phi8*/	7,46,4,5,47,1,8,64,2,6,64,3,9,127,1,1,134,2,1,135,0,11,
/* out0173_em-eta13-phi8*/	6,46,1,2,46,2,7,47,0,10,47,1,6,127,1,10,127,2,1,
/* out0174_em-eta14-phi8*/	6,46,2,8,46,3,4,47,3,2,47,4,6,127,0,4,127,2,4,
/* out0175_em-eta15-phi8*/	9,27,2,1,29,1,3,46,3,4,47,3,8,119,1,3,119,2,1,120,0,1,127,0,2,127,2,1,
/* out0176_em-eta16-phi8*/	4,28,1,10,28,2,1,29,1,4,119,2,6,
/* out0177_em-eta17-phi8*/	5,28,0,4,28,1,5,28,2,3,112,1,1,119,2,4,
/* out0178_em-eta18-phi8*/	3,28,0,4,28,3,6,112,1,4,
/* out0179_em-eta19-phi8*/	2,11,0,3,28,3,4,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	3,134,2,7,135,0,3,135,1,3,
/* out0183_em-eta3-phi9*/	6,127,0,3,127,1,16,127,2,3,134,0,7,134,2,6,135,0,10,
/* out0184_em-eta4-phi9*/	6,116,1,1,116,2,1,117,0,2,117,1,9,127,0,6,127,2,12,
/* out0185_em-eta5-phi9*/	6,104,2,5,105,1,1,116,2,1,117,0,14,117,1,1,117,2,5,
/* out0186_em-eta6-phi9*/	5,92,1,1,104,0,3,104,2,9,105,0,9,105,1,1,
/* out0187_em-eta7-phi9*/	4,92,0,1,92,1,5,92,2,11,105,0,1,
/* out0188_em-eta8-phi9*/	3,80,1,4,92,0,8,92,2,2,
/* out0189_em-eta9-phi9*/	3,80,0,3,80,1,9,80,2,1,
/* out0190_em-eta10-phi9*/	4,63,5,7,64,5,1,66,1,3,80,0,8,
/* out0191_em-eta11-phi9*/	8,64,2,4,64,5,10,65,0,4,65,1,15,66,1,2,135,1,7,135,2,6,136,0,1,
/* out0192_em-eta12-phi9*/	8,46,4,10,46,5,1,64,2,3,65,0,12,65,3,3,128,1,1,135,0,2,135,2,9,
/* out0193_em-eta13-phi9*/	10,46,4,1,46,5,12,47,0,6,47,4,3,47,5,3,127,1,1,127,2,4,128,0,4,128,1,1,135,0,1,
/* out0194_em-eta14-phi9*/	7,47,2,5,47,3,3,47,4,7,47,5,5,120,1,2,127,2,6,128,0,1,
/* out0195_em-eta15-phi9*/	6,28,4,5,29,1,3,47,2,6,47,3,3,120,0,2,120,1,5,
/* out0196_em-eta16-phi9*/	5,28,2,1,28,4,1,29,0,6,29,1,6,120,0,6,
/* out0197_em-eta17-phi9*/	6,28,2,8,29,0,3,29,4,2,112,1,2,112,2,3,120,0,1,
/* out0198_em-eta18-phi9*/	6,28,2,3,28,3,3,29,3,2,29,4,2,112,1,5,112,2,1,
/* out0199_em-eta19-phi9*/	2,28,3,3,29,3,5,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	2,135,1,10,135,2,1,
/* out0203_em-eta3-phi10*/	7,127,2,1,128,1,9,128,2,4,135,0,3,135,1,3,135,2,15,136,0,7,
/* out0204_em-eta4-phi10*/	5,117,1,5,118,1,2,128,0,14,128,1,7,128,2,3,
/* out0205_em-eta5-phi10*/	5,105,1,4,117,1,1,117,2,11,118,0,10,118,1,1,
/* out0206_em-eta6-phi10*/	3,105,0,4,105,1,10,105,2,8,
/* out0207_em-eta7-phi10*/	4,92,2,2,93,1,10,105,0,2,105,2,5,
/* out0208_em-eta8-phi10*/	4,80,2,2,92,2,1,93,0,7,93,1,4,
/* out0209_em-eta9-phi10*/	3,80,2,11,81,1,1,93,0,1,
/* out0210_em-eta10-phi10*/	5,65,4,12,66,1,5,80,0,4,80,2,2,81,1,1,
/* out0211_em-eta11-phi10*/	9,65,1,1,65,2,9,65,4,1,65,5,1,66,0,13,66,1,6,66,4,3,136,0,11,136,2,2,
/* out0212_em-eta12-phi10*/	8,65,2,7,65,3,10,66,3,6,66,4,5,128,1,9,135,2,1,136,0,1,136,2,4,
/* out0213_em-eta13-phi10*/	9,46,5,3,47,5,5,48,1,5,49,1,4,65,3,3,66,3,4,128,0,5,128,1,3,128,2,2,
/* out0214_em-eta14-phi10*/	6,47,2,4,47,5,3,48,0,7,48,1,7,120,1,4,128,0,5,
/* out0215_em-eta15-phi10*/	5,28,4,8,47,2,1,48,0,8,120,1,5,120,2,3,
/* out0216_em-eta16-phi10*/	5,28,4,2,28,5,8,29,0,4,120,0,4,120,2,2,
/* out0217_em-eta17-phi10*/	5,29,0,3,29,4,8,29,5,1,112,2,4,120,0,2,
/* out0218_em-eta18-phi10*/	5,29,2,2,29,3,4,29,4,4,112,1,2,112,2,4,
/* out0219_em-eta19-phi10*/	3,29,2,1,29,3,5,112,1,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	4,128,2,3,129,1,7,136,0,9,136,2,16,
/* out0224_em-eta4-phi11*/	5,118,1,7,128,0,2,128,2,6,129,0,8,129,1,9,
/* out0225_em-eta5-phi11*/	4,106,1,1,118,0,5,118,1,6,118,2,15,
/* out0226_em-eta6-phi11*/	5,105,2,3,106,0,10,106,1,7,118,0,1,118,2,1,
/* out0227_em-eta7-phi11*/	3,93,1,2,93,2,10,106,0,6,
/* out0228_em-eta8-phi11*/	3,81,1,1,93,0,8,93,2,6,
/* out0229_em-eta9-phi11*/	1,81,1,12,
/* out0230_em-eta10-phi11*/	4,65,4,3,65,5,3,81,0,8,81,1,1,
/* out0231_em-eta11-phi11*/	7,65,5,12,66,0,3,66,4,5,66,5,14,129,1,2,136,0,3,136,2,7,
/* out0232_em-eta12-phi11*/	10,48,4,3,66,2,16,66,3,5,66,4,3,66,5,2,128,1,2,128,2,3,129,0,3,129,1,2,136,2,3,
/* out0233_em-eta13-phi11*/	8,48,1,1,48,4,5,49,0,5,49,1,12,66,3,1,121,1,1,128,2,9,129,0,1,
/* out0234_em-eta14-phi11*/	8,48,1,3,48,2,14,49,0,3,120,2,1,121,0,2,121,1,3,128,0,1,128,2,2,
/* out0235_em-eta15-phi11*/	5,48,0,1,48,2,2,48,3,13,120,2,5,121,0,2,
/* out0236_em-eta16-phi11*/	5,28,5,8,29,5,4,48,3,3,113,1,2,120,2,4,
/* out0237_em-eta17-phi11*/	6,29,2,1,29,5,11,112,2,1,113,0,2,113,1,2,120,2,1,
/* out0238_em-eta18-phi11*/	3,29,2,10,112,2,3,113,0,2,
/* out0239_em-eta19-phi11*/	2,29,2,2,112,1,1,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	4,129,2,7,130,1,3,137,1,9,137,2,16,
/* out0244_em-eta4-phi12*/	6,119,1,4,119,2,3,129,0,8,129,2,9,130,0,2,130,1,6,
/* out0245_em-eta5-phi12*/	4,106,1,1,119,0,11,119,1,12,119,2,3,
/* out0246_em-eta6-phi12*/	4,106,1,7,106,2,10,107,0,3,119,0,1,
/* out0247_em-eta7-phi12*/	3,94,0,2,94,1,10,106,2,6,
/* out0248_em-eta8-phi12*/	2,81,2,1,94,0,13,
/* out0249_em-eta9-phi12*/	2,81,2,12,94,0,1,
/* out0250_em-eta10-phi12*/	4,67,4,1,67,5,5,81,0,8,81,2,1,
/* out0251_em-eta11-phi12*/	6,67,4,15,67,5,5,68,0,7,68,1,7,129,1,8,129,2,1,
/* out0252_em-eta12-phi12*/	8,48,4,3,67,1,13,67,2,2,68,0,2,68,1,9,129,0,6,129,1,4,129,2,3,
/* out0253_em-eta13-phi12*/	7,48,4,5,48,5,12,49,0,5,49,5,1,67,0,1,121,1,6,129,0,5,
/* out0254_em-eta14-phi12*/	6,49,0,3,49,4,14,49,5,3,121,0,3,121,1,5,121,2,1,
/* out0255_em-eta15-phi12*/	4,49,2,1,49,3,13,49,4,2,121,0,7,
/* out0256_em-eta16-phi12*/	3,30,4,11,49,3,3,113,1,6,
/* out0257_em-eta17-phi12*/	4,30,4,5,31,1,7,113,0,3,113,1,3,
/* out0258_em-eta18-phi12*/	3,30,1,3,31,1,7,113,0,4,
/* out0259_em-eta19-phi12*/	2,30,1,2,113,0,1,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	2,138,0,2,138,1,5,
/* out0263_em-eta3-phi13*/	7,130,1,4,130,2,9,131,0,1,137,1,7,138,0,14,138,1,3,138,2,12,
/* out0264_em-eta4-phi13*/	5,119,2,2,120,1,6,130,0,14,130,1,3,130,2,7,
/* out0265_em-eta5-phi13*/	5,107,1,4,119,0,4,119,2,8,120,0,3,120,1,8,
/* out0266_em-eta6-phi13*/	3,107,0,8,107,1,10,107,2,4,
/* out0267_em-eta7-phi13*/	5,94,1,6,94,2,4,95,0,1,107,0,5,107,2,2,
/* out0268_em-eta8-phi13*/	3,82,1,2,94,2,12,95,0,1,
/* out0269_em-eta9-phi13*/	2,81,2,1,82,1,11,
/* out0270_em-eta10-phi13*/	6,67,5,4,68,2,2,68,5,11,81,2,1,82,0,4,82,1,2,
/* out0271_em-eta11-phi13*/	9,67,2,2,67,5,2,68,0,7,68,2,2,68,3,1,68,4,16,68,5,5,129,2,3,130,0,9,
/* out0272_em-eta12-phi13*/	7,67,0,8,67,1,3,67,2,12,67,3,6,122,1,3,129,2,8,130,0,1,
/* out0273_em-eta13-phi13*/	10,48,5,4,49,5,5,50,4,9,67,0,7,121,1,1,121,2,2,122,0,3,122,1,2,129,0,1,129,2,1,
/* out0274_em-eta14-phi13*/	5,49,2,7,49,5,7,50,4,1,51,1,5,121,2,9,
/* out0275_em-eta15-phi13*/	7,30,5,7,31,5,2,49,2,8,51,1,1,114,1,1,121,0,2,121,2,3,
/* out0276_em-eta16-phi13*/	4,30,5,9,31,0,4,113,1,3,113,2,4,
/* out0277_em-eta17-phi13*/	4,30,2,1,31,0,10,31,1,1,113,2,5,
/* out0278_em-eta18-phi13*/	6,30,1,6,30,2,3,31,0,1,31,1,1,113,0,3,113,2,1,
/* out0279_em-eta19-phi13*/	3,30,0,3,30,1,4,113,0,1,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	2,138,1,4,139,0,7,
/* out0283_em-eta3-phi14*/	7,131,0,3,131,1,16,131,2,3,138,1,4,138,2,4,139,0,6,139,2,7,
/* out0284_em-eta4-phi14*/	5,120,1,1,120,2,10,121,1,3,131,0,12,131,2,6,
/* out0285_em-eta5-phi14*/	6,107,1,1,108,1,5,120,0,13,120,1,1,120,2,6,121,1,1,
/* out0286_em-eta6-phi14*/	5,95,1,1,107,1,1,107,2,9,108,0,3,108,1,9,
/* out0287_em-eta7-phi14*/	4,95,0,4,95,1,12,95,2,1,107,2,1,
/* out0288_em-eta8-phi14*/	3,82,2,4,95,0,10,95,2,1,
/* out0289_em-eta9-phi14*/	3,82,0,3,82,1,1,82,2,9,
/* out0290_em-eta10-phi14*/	3,68,2,3,69,4,7,82,0,8,
/* out0291_em-eta11-phi14*/	6,68,2,9,68,3,11,69,4,7,70,1,7,130,0,6,130,2,12,
/* out0292_em-eta12-phi14*/	9,50,5,8,51,5,2,67,3,10,68,3,4,69,1,1,70,1,2,122,1,9,122,2,2,130,2,2,
/* out0293_em-eta13-phi14*/	7,50,4,6,50,5,8,51,0,9,51,1,1,122,0,8,122,1,2,122,2,2,
/* out0294_em-eta14-phi14*/	7,50,1,5,50,2,3,51,0,5,51,1,9,114,1,5,121,2,1,122,0,3,
/* out0295_em-eta15-phi14*/	5,31,2,1,31,5,7,50,1,8,114,0,2,114,1,6,
/* out0296_em-eta16-phi14*/	4,31,4,7,31,5,7,113,2,1,114,0,5,
/* out0297_em-eta17-phi14*/	5,30,2,5,31,0,1,31,4,6,107,1,1,113,2,3,
/* out0298_em-eta18-phi14*/	6,30,0,1,30,1,1,30,2,6,30,3,2,107,1,2,113,2,2,
/* out0299_em-eta19-phi14*/	2,30,0,8,107,1,1,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	1,139,0,1,
/* out0303_em-eta3-phi15*/	6,131,2,4,132,0,11,132,1,14,132,2,2,139,0,2,139,2,9,
/* out0304_em-eta4-phi15*/	5,121,0,2,121,1,10,121,2,12,131,2,3,132,0,5,
/* out0305_em-eta5-phi15*/	5,108,1,1,108,2,10,109,1,2,121,0,12,121,1,2,
/* out0306_em-eta6-phi15*/	4,96,1,2,108,0,13,108,1,1,108,2,6,
/* out0307_em-eta7-phi15*/	3,95,1,3,95,2,8,96,1,6,
/* out0308_em-eta8-phi15*/	3,83,1,8,83,2,1,95,2,6,
/* out0309_em-eta9-phi15*/	3,82,2,3,83,0,3,83,1,7,
/* out0310_em-eta10-phi15*/	6,69,4,1,69,5,16,70,0,4,70,4,5,70,5,12,82,0,1,
/* out0311_em-eta11-phi15*/	10,69,1,4,69,2,9,69,4,1,70,0,12,70,1,7,70,4,2,123,0,16,123,1,4,123,2,2,130,2,2,
/* out0312_em-eta12-phi15*/	7,51,2,4,51,5,10,69,0,4,69,1,11,115,1,1,122,2,6,123,2,8,
/* out0313_em-eta13-phi15*/	8,51,0,2,51,2,2,51,3,1,51,4,15,51,5,4,115,1,3,122,0,1,122,2,6,
/* out0314_em-eta14-phi15*/	9,50,0,1,50,1,2,50,2,13,50,3,3,51,4,1,114,1,3,114,2,4,115,0,1,122,0,1,
/* out0315_em-eta15-phi15*/	7,31,2,4,32,1,1,50,0,12,50,1,1,114,0,2,114,1,1,114,2,5,
/* out0316_em-eta16-phi15*/	4,31,2,10,31,3,3,31,4,1,114,0,6,
/* out0317_em-eta17-phi15*/	6,30,2,1,30,3,1,31,3,8,31,4,2,107,1,1,107,2,4,
/* out0318_em-eta18-phi15*/	2,30,3,10,107,1,4,
/* out0319_em-eta19-phi15*/	3,13,4,3,30,0,4,107,1,2,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	2,133,0,3,133,2,1,
/* out0323_em-eta3-phi16*/	6,122,1,1,122,2,3,132,1,2,132,2,12,133,0,13,133,2,12,
/* out0324_em-eta4-phi16*/	5,121,2,4,122,0,8,122,1,15,122,2,4,132,2,2,
/* out0325_em-eta5-phi16*/	4,109,0,3,109,1,12,109,2,9,121,0,2,
/* out0326_em-eta6-phi16*/	4,96,1,3,96,2,8,109,0,7,109,1,2,
/* out0327_em-eta7-phi16*/	3,96,0,10,96,1,5,96,2,3,
/* out0328_em-eta8-phi16*/	3,83,1,1,83,2,12,96,0,3,
/* out0329_em-eta9-phi16*/	2,83,0,10,83,2,1,
/* out0330_em-eta10-phi16*/	6,70,2,16,70,3,6,70,4,4,70,5,4,71,1,2,83,0,1,
/* out0331_em-eta11-phi16*/	5,69,2,7,69,3,14,70,3,8,70,4,5,123,1,10,
/* out0332_em-eta12-phi16*/	8,51,2,4,52,1,4,53,1,8,69,0,12,115,1,5,115,2,1,123,1,2,123,2,6,
/* out0333_em-eta13-phi16*/	7,51,2,6,51,3,11,52,0,3,52,1,5,115,0,2,115,1,7,115,2,1,
/* out0334_em-eta14-phi16*/	5,32,4,3,50,3,13,51,3,4,114,2,1,115,0,7,
/* out0335_em-eta15-phi16*/	6,32,1,1,32,4,1,33,1,13,50,0,3,108,1,3,114,2,5,
/* out0336_em-eta16-phi16*/	8,31,2,1,32,0,1,32,1,12,107,2,2,108,0,1,108,1,2,114,0,1,114,2,1,
/* out0337_em-eta17-phi16*/	3,31,3,5,32,0,6,107,2,6,
/* out0338_em-eta18-phi16*/	6,13,5,10,14,5,1,30,3,3,107,0,2,107,1,2,107,2,1,
/* out0339_em-eta19-phi16*/	3,13,4,8,13,5,1,107,1,2,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	2,122,2,2,133,2,3,
/* out0344_em-eta4-phi17*/	4,110,1,10,122,0,8,122,2,7,123,2,5,
/* out0345_em-eta5-phi17*/	5,97,1,3,109,0,3,109,2,7,110,0,12,110,1,2,
/* out0346_em-eta6-phi17*/	4,96,2,2,97,0,8,97,1,9,109,0,3,
/* out0347_em-eta7-phi17*/	5,84,1,5,84,2,4,96,0,3,96,2,3,97,0,4,
/* out0348_em-eta8-phi17*/	3,83,2,1,84,0,3,84,1,11,
/* out0349_em-eta9-phi17*/	5,71,1,5,71,2,4,83,0,2,83,2,1,84,0,1,
/* out0350_em-eta10-phi17*/	2,71,0,2,71,1,8,
/* out0351_em-eta11-phi17*/	8,52,4,14,52,5,3,69,3,2,70,3,2,71,0,2,71,1,1,116,0,12,116,1,5,
/* out0352_em-eta12-phi17*/	9,52,1,2,52,2,5,52,4,2,52,5,1,53,0,12,53,1,8,115,2,3,116,0,4,116,2,8,
/* out0353_em-eta13-phi17*/	6,52,0,8,52,1,5,52,2,7,52,3,3,115,0,1,115,2,10,
/* out0354_em-eta14-phi17*/	7,32,4,11,32,5,3,52,0,5,52,3,1,108,1,3,115,0,5,115,2,1,
/* out0355_em-eta15-phi17*/	5,32,4,1,32,5,1,33,0,12,33,1,3,108,1,7,
/* out0356_em-eta16-phi17*/	4,32,1,2,32,2,12,108,0,5,108,1,1,
/* out0357_em-eta17-phi17*/	5,32,0,8,32,3,4,107,0,1,107,2,3,108,0,2,
/* out0358_em-eta18-phi17*/	6,13,5,3,14,0,2,14,4,3,14,5,11,32,0,1,107,0,10,
/* out0359_em-eta19-phi17*/	7,13,4,5,13,5,2,14,0,10,14,1,2,14,4,1,107,0,3,107,1,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	2,124,0,2,124,1,4,
/* out0363_em-eta3-phi18*/	7,111,1,1,111,2,1,123,1,12,123,2,5,124,0,14,124,1,2,124,2,3,
/* out0364_em-eta4-phi18*/	7,110,1,4,110,2,6,111,0,1,111,1,14,111,2,1,123,1,4,123,2,6,
/* out0365_em-eta5-phi18*/	6,97,1,2,97,2,1,98,1,9,98,2,1,110,0,4,110,2,10,
/* out0366_em-eta6-phi18*/	5,85,1,2,97,0,1,97,1,2,97,2,14,98,1,3,
/* out0367_em-eta7-phi18*/	4,84,2,8,85,1,6,97,0,3,97,2,1,
/* out0368_em-eta8-phi18*/	3,72,1,1,84,0,10,84,2,4,
/* out0369_em-eta9-phi18*/	3,71,2,8,72,1,2,84,0,2,
/* out0370_em-eta10-phi18*/	2,71,0,8,71,2,3,
/* out0371_em-eta11-phi18*/	6,52,5,11,53,5,6,54,4,4,71,0,3,110,0,1,116,1,9,
/* out0372_em-eta12-phi18*/	9,52,5,1,53,0,4,53,2,1,53,3,1,53,4,12,53,5,9,109,1,3,116,1,2,116,2,8,
/* out0373_em-eta13-phi18*/	6,52,2,4,52,3,7,53,3,10,53,4,4,109,0,1,109,1,10,
/* out0374_em-eta14-phi18*/	7,32,5,11,33,5,4,52,3,5,53,3,1,108,2,3,109,0,5,109,1,1,
/* out0375_em-eta15-phi18*/	5,32,5,1,33,0,4,33,4,8,33,5,4,108,2,7,
/* out0376_em-eta16-phi18*/	5,32,2,4,33,3,2,33,4,8,108,0,5,108,2,1,
/* out0377_em-eta17-phi18*/	5,32,3,10,33,3,2,103,1,1,103,2,3,108,0,2,
/* out0378_em-eta18-phi18*/	6,14,2,8,14,3,1,14,4,2,14,5,4,32,3,1,103,1,4,
/* out0379_em-eta19-phi18*/	6,13,1,4,13,3,4,14,0,4,14,1,8,14,4,9,103,1,2,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	1,124,1,2,
/* out0383_em-eta3-phi19*/	5,111,2,5,112,1,12,112,2,2,124,1,8,124,2,13,
/* out0384_em-eta4-phi19*/	5,99,1,4,111,0,15,111,1,1,111,2,9,112,1,2,
/* out0385_em-eta5-phi19*/	4,98,0,6,98,1,3,98,2,15,99,0,2,
/* out0386_em-eta6-phi19*/	4,85,1,1,85,2,10,98,0,9,98,1,1,
/* out0387_em-eta7-phi19*/	3,85,0,9,85,1,7,85,2,3,
/* out0388_em-eta8-phi19*/	3,72,1,5,72,2,8,85,0,2,
/* out0389_em-eta9-phi19*/	2,72,0,5,72,1,8,
/* out0390_em-eta10-phi19*/	8,54,4,1,54,5,13,55,0,2,55,4,2,55,5,12,71,0,1,71,2,1,72,0,1,
/* out0391_em-eta11-phi19*/	7,54,4,11,54,5,3,55,0,12,55,1,8,110,0,12,110,1,5,110,2,1,
/* out0392_em-eta12-phi19*/	10,34,5,2,35,5,2,53,2,12,53,5,1,54,1,4,55,1,8,109,1,1,109,2,5,110,0,3,110,2,7,
/* out0393_em-eta13-phi19*/	7,34,4,5,34,5,12,53,2,3,53,3,4,109,0,2,109,1,1,109,2,7,
/* out0394_em-eta14-phi19*/	6,33,5,3,34,4,11,35,0,1,35,1,5,104,1,1,109,0,7,
/* out0395_em-eta15-phi19*/	5,33,2,9,33,5,5,35,1,3,104,1,5,108,2,3,
/* out0396_em-eta16-phi19*/	8,15,5,1,33,2,6,33,3,6,103,2,2,104,0,1,104,1,1,108,0,1,108,2,2,
/* out0397_em-eta17-phi19*/	4,15,4,5,32,3,1,33,3,6,103,2,6,
/* out0398_em-eta18-phi19*/	5,14,2,8,14,3,2,15,4,3,103,1,3,103,2,1,
/* out0399_em-eta19-phi19*/	6,13,1,10,13,3,10,14,1,5,14,3,9,14,4,1,103,1,2,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	1,113,2,1,
/* out0403_em-eta3-phi20*/	6,100,1,4,112,0,11,112,1,2,112,2,14,113,0,9,113,2,2,
/* out0404_em-eta4-phi20*/	5,99,0,2,99,1,12,99,2,10,100,1,3,112,0,5,
/* out0405_em-eta5-phi20*/	5,86,1,10,86,2,1,98,0,1,99,0,12,99,2,2,
/* out0406_em-eta6-phi20*/	4,85,2,2,86,0,13,86,1,6,86,2,1,
/* out0407_em-eta7-phi20*/	4,73,1,8,73,2,3,85,0,5,85,2,1,
/* out0408_em-eta8-phi20*/	3,72,0,1,72,2,8,73,1,6,
/* out0409_em-eta9-phi20*/	2,56,1,3,72,0,9,
/* out0410_em-eta10-phi20*/	5,55,2,16,55,3,8,55,4,9,55,5,4,56,0,1,
/* out0411_em-eta11-phi20*/	10,54,0,3,54,1,3,54,2,16,54,3,5,55,0,2,55,3,1,55,4,5,106,0,2,110,1,11,110,2,1,
/* out0412_em-eta12-phi20*/	7,35,2,5,35,5,8,54,0,6,54,1,9,105,1,6,109,2,1,110,2,7,
/* out0413_em-eta13-phi20*/	7,34,5,2,35,0,7,35,4,10,35,5,6,105,0,1,105,1,6,109,2,3,
/* out0414_em-eta14-phi20*/	8,34,1,2,34,2,6,35,0,8,35,1,4,104,1,4,104,2,3,105,0,1,109,0,1,
/* out0415_em-eta15-phi20*/	7,16,5,3,33,2,1,34,1,8,35,1,4,104,0,2,104,1,5,104,2,1,
/* out0416_em-eta16-phi20*/	4,15,5,10,16,0,1,16,5,4,104,0,6,
/* out0417_em-eta17-phi20*/	5,15,4,4,15,5,5,16,0,3,103,0,2,103,2,4,
/* out0418_em-eta18-phi20*/	4,15,4,4,16,1,6,103,0,5,103,1,2,
/* out0419_em-eta19-phi20*/	6,13,1,2,13,3,2,14,1,1,14,3,4,16,1,4,103,1,1,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	3,101,0,3,101,1,3,113,2,7,
/* out0423_em-eta3-phi21*/	6,100,0,3,100,1,3,100,2,16,101,0,10,113,0,7,113,2,6,
/* out0424_em-eta4-phi21*/	5,87,1,10,87,2,1,99,2,3,100,0,12,100,1,6,
/* out0425_em-eta5-phi21*/	6,74,2,1,86,2,5,87,0,13,87,1,6,87,2,1,99,2,1,
/* out0426_em-eta6-phi21*/	5,73,2,1,74,1,9,74,2,1,86,0,3,86,2,9,
/* out0427_em-eta7-phi21*/	4,73,0,4,73,1,1,73,2,12,74,1,1,
/* out0428_em-eta8-phi21*/	3,56,1,4,73,0,10,73,1,1,
/* out0429_em-eta9-phi21*/	3,56,0,3,56,1,9,56,2,1,
/* out0430_em-eta10-phi21*/	4,36,4,3,54,3,1,55,3,7,56,0,8,
/* out0431_em-eta11-phi21*/	6,36,4,9,37,1,11,54,0,4,54,3,10,106,0,12,106,2,6,
/* out0432_em-eta12-phi21*/	8,35,2,10,35,3,1,36,1,10,37,1,4,54,0,3,105,1,2,105,2,9,106,2,2,
/* out0433_em-eta13-phi21*/	8,34,2,3,34,3,3,35,2,1,35,3,12,35,4,6,105,0,8,105,1,2,105,2,2,
/* out0434_em-eta14-phi21*/	7,34,0,5,34,1,3,34,2,7,34,3,5,101,1,1,104,2,5,105,0,3,
/* out0435_em-eta15-phi21*/	6,16,2,5,16,5,3,34,0,6,34,1,3,104,0,2,104,2,6,
/* out0436_em-eta16-phi21*/	6,16,0,1,16,2,1,16,4,6,16,5,6,100,1,1,104,0,5,
/* out0437_em-eta17-phi21*/	5,15,2,2,16,0,8,16,4,3,100,1,3,103,0,3,
/* out0438_em-eta18-phi21*/	6,15,1,2,15,2,2,16,0,3,16,1,3,100,1,2,103,0,6,
/* out0439_em-eta19-phi21*/	4,15,1,5,16,1,3,100,0,1,103,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	2,101,1,10,101,2,1,
/* out0443_em-eta3-phi22*/	7,88,1,9,88,2,4,89,0,7,100,0,1,101,0,3,101,1,3,101,2,15,
/* out0444_em-eta4-phi22*/	5,75,1,2,87,2,6,88,0,14,88,1,7,88,2,3,
/* out0445_em-eta5-phi22*/	5,74,2,4,75,0,4,75,1,8,87,0,3,87,2,8,
/* out0446_em-eta6-phi22*/	3,74,0,8,74,1,4,74,2,10,
/* out0447_em-eta7-phi22*/	5,57,1,4,57,2,6,73,0,1,74,0,5,74,1,2,
/* out0448_em-eta8-phi22*/	3,56,2,2,57,1,12,73,0,1,
/* out0449_em-eta9-phi22*/	2,38,1,1,56,2,11,
/* out0450_em-eta10-phi22*/	7,36,4,2,36,5,11,37,5,4,38,0,6,38,1,1,56,0,4,56,2,2,
/* out0451_em-eta11-phi22*/	11,36,2,2,36,4,2,36,5,5,37,0,16,37,1,1,37,4,7,37,5,2,102,1,3,102,2,3,106,0,2,106,2,7,
/* out0452_em-eta12-phi22*/	8,36,0,8,36,1,6,36,2,12,36,3,3,102,0,3,102,1,8,105,2,3,106,2,1,
/* out0453_em-eta13-phi22*/	11,17,5,5,18,5,4,34,3,5,35,3,3,36,0,7,101,1,2,101,2,2,102,0,1,102,1,1,105,0,3,105,2,2,
/* out0454_em-eta14-phi22*/	6,17,4,7,17,5,7,34,0,4,34,3,3,101,1,9,101,2,2,
/* out0455_em-eta15-phi22*/	7,16,2,8,17,4,8,34,0,1,100,2,1,101,0,5,101,1,3,104,2,1,
/* out0456_em-eta16-phi22*/	5,16,2,2,16,3,8,16,4,4,100,1,4,100,2,3,
/* out0457_em-eta17-phi22*/	6,15,2,8,15,3,1,16,4,3,100,0,1,100,1,5,100,2,1,
/* out0458_em-eta18-phi22*/	5,15,0,2,15,1,4,15,2,4,100,0,4,100,1,1,
/* out0459_em-eta19-phi22*/	3,15,0,1,15,1,5,100,0,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	4,76,1,7,88,2,3,89,0,9,89,2,16,
/* out0464_em-eta4-phi23*/	6,75,1,3,75,2,4,76,0,16,76,1,9,88,0,2,88,2,6,
/* out0465_em-eta5-phi23*/	4,58,2,9,75,0,11,75,1,3,75,2,12,
/* out0466_em-eta6-phi23*/	4,58,1,10,58,2,7,74,0,3,75,0,1,
/* out0467_em-eta7-phi23*/	3,57,0,2,57,2,10,58,1,6,
/* out0468_em-eta8-phi23*/	3,38,1,1,38,2,15,57,0,13,
/* out0469_em-eta9-phi23*/	4,38,0,1,38,1,12,38,2,1,57,0,1,
/* out0470_em-eta10-phi23*/	4,37,2,1,37,5,5,38,0,8,38,1,1,
/* out0471_em-eta11-phi23*/	7,37,2,15,37,3,7,37,4,7,37,5,5,38,0,1,102,1,1,102,2,9,
/* out0472_em-eta12-phi23*/	8,18,2,3,36,2,2,36,3,13,37,3,9,37,4,2,102,0,7,102,1,3,102,2,4,
/* out0473_em-eta13-phi23*/	7,17,5,1,18,2,13,18,4,13,18,5,12,36,0,1,101,2,6,102,0,5,
/* out0474_em-eta14-phi23*/	6,17,5,3,18,0,14,18,4,3,101,0,3,101,1,1,101,2,6,
/* out0475_em-eta15-phi23*/	5,17,4,1,18,0,2,18,1,13,100,2,1,101,0,8,
/* out0476_em-eta16-phi23*/	5,15,3,4,16,3,8,17,1,16,18,1,3,100,2,7,
/* out0477_em-eta17-phi23*/	4,15,0,1,15,3,11,100,0,3,100,2,3,
/* out0478_em-eta18-phi23*/	2,15,0,10,100,0,5,
/* out0479_em-eta19-phi23*/	2,15,0,2,100,0,1
};