parameter integer matrixH [0:5042] = {
/* num inputs = 152(in0-in151) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1520 */

/* out0000_em-eta0-phi0*/	1,107,0,4,
/* out0001_em-eta1-phi0*/	2,106,0,6,107,0,12,
/* out0002_em-eta2-phi0*/	2,106,0,10,106,1,8,
/* out0003_em-eta3-phi0*/	2,105,0,9,106,1,8,
/* out0004_em-eta4-phi0*/	2,105,0,7,105,1,10,
/* out0005_em-eta5-phi0*/	2,104,0,11,105,1,6,
/* out0006_em-eta6-phi0*/	2,104,0,5,104,1,16,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	5,47,0,13,47,1,12,47,2,2,99,1,3,99,2,13,
/* out0010_em-eta10-phi0*/	6,46,0,1,46,1,4,47,0,3,47,2,9,98,0,9,98,1,3,
/* out0011_em-eta11-phi0*/	5,46,0,6,46,1,6,46,2,2,98,0,7,98,2,2,
/* out0012_em-eta12-phi0*/	6,45,0,6,45,1,2,46,0,9,46,2,7,97,0,8,97,1,1,
/* out0013_em-eta13-phi0*/	3,45,0,5,45,1,5,97,0,6,
/* out0014_em-eta14-phi0*/	3,45,0,4,45,2,5,96,0,3,
/* out0015_em-eta15-phi0*/	5,44,0,7,44,1,4,45,0,1,45,2,2,96,0,6,
/* out0016_em-eta16-phi0*/	3,44,0,5,44,1,1,96,0,2,
/* out0017_em-eta17-phi0*/	3,44,0,3,44,2,2,95,0,2,
/* out0018_em-eta18-phi0*/	3,44,0,1,44,2,1,95,0,3,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	1,107,1,4,
/* out0021_em-eta1-phi1*/	2,106,3,6,107,1,12,
/* out0022_em-eta2-phi1*/	2,106,2,8,106,3,10,
/* out0023_em-eta3-phi1*/	2,105,3,9,106,2,8,
/* out0024_em-eta4-phi1*/	2,105,2,10,105,3,7,
/* out0025_em-eta5-phi1*/	2,104,3,11,105,2,6,
/* out0026_em-eta6-phi1*/	2,104,2,16,104,3,5,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	1,43,2,2,
/* out0029_em-eta9-phi1*/	9,42,0,1,42,1,2,43,1,4,43,2,11,47,1,4,47,2,2,93,0,5,99,1,13,99,2,3,
/* out0030_em-eta10-phi1*/	7,42,0,11,42,1,1,46,1,1,47,2,3,93,0,2,98,1,12,98,2,2,
/* out0031_em-eta11-phi1*/	8,41,0,1,42,0,3,42,2,1,46,1,5,46,2,3,91,0,1,97,1,2,98,2,11,
/* out0032_em-eta12-phi1*/	6,41,0,6,45,1,2,46,2,4,97,0,1,97,1,10,97,2,1,
/* out0033_em-eta13-phi1*/	5,41,0,2,45,1,7,45,2,1,97,0,1,97,2,9,
/* out0034_em-eta14-phi1*/	5,40,0,1,45,2,7,96,0,1,96,1,7,97,2,1,
/* out0035_em-eta15-phi1*/	6,40,0,1,44,1,5,45,2,1,96,0,3,96,1,1,96,2,2,
/* out0036_em-eta16-phi1*/	5,44,1,4,44,2,2,95,1,1,96,0,1,96,2,4,
/* out0037_em-eta17-phi1*/	3,44,2,5,95,0,4,95,1,3,
/* out0038_em-eta18-phi1*/	2,44,2,2,95,0,3,
/* out0039_em-eta19-phi1*/	0,
/* out0040_em-eta0-phi2*/	1,111,0,4,
/* out0041_em-eta1-phi2*/	2,110,0,6,111,0,12,
/* out0042_em-eta2-phi2*/	2,110,0,10,110,1,8,
/* out0043_em-eta3-phi2*/	2,109,0,9,110,1,8,
/* out0044_em-eta4-phi2*/	2,109,0,7,109,1,10,
/* out0045_em-eta5-phi2*/	2,108,0,11,109,1,6,
/* out0046_em-eta6-phi2*/	2,108,0,5,108,1,16,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	5,37,0,1,37,2,1,43,1,2,43,2,3,93,1,1,
/* out0049_em-eta9-phi2*/	6,37,2,9,42,1,5,43,1,10,93,0,5,93,1,13,93,2,3,
/* out0050_em-eta10-phi2*/	9,42,0,1,42,1,8,42,2,8,91,0,1,91,1,4,93,0,4,93,2,8,98,1,1,98,2,1,
/* out0051_em-eta11-phi2*/	5,41,1,7,42,2,6,91,0,11,91,1,3,91,2,1,
/* out0052_em-eta12-phi2*/	9,41,0,5,41,1,4,41,2,3,90,0,1,90,1,1,91,0,3,91,2,2,97,1,3,97,2,2,
/* out0053_em-eta13-phi2*/	5,40,1,2,41,0,2,41,2,4,90,0,6,97,2,3,
/* out0054_em-eta14-phi2*/	4,40,0,6,40,1,2,90,0,3,96,1,6,
/* out0055_em-eta15-phi2*/	3,40,0,6,96,1,2,96,2,5,
/* out0056_em-eta16-phi2*/	7,39,1,1,40,0,1,44,1,2,44,2,2,89,0,1,95,1,2,96,2,4,
/* out0057_em-eta17-phi2*/	3,39,1,2,44,2,2,95,1,6,
/* out0058_em-eta18-phi2*/	3,39,0,1,39,1,1,95,0,3,
/* out0059_em-eta19-phi2*/	0,
/* out0060_em-eta0-phi3*/	1,111,1,4,
/* out0061_em-eta1-phi3*/	2,110,3,6,111,1,12,
/* out0062_em-eta2-phi3*/	2,110,2,8,110,3,10,
/* out0063_em-eta3-phi3*/	2,109,3,9,110,2,8,
/* out0064_em-eta4-phi3*/	2,109,2,10,109,3,7,
/* out0065_em-eta5-phi3*/	2,108,3,11,109,2,6,
/* out0066_em-eta6-phi3*/	2,108,2,16,108,3,5,
/* out0067_em-eta7-phi3*/	0,
/* out0068_em-eta8-phi3*/	1,37,0,5,
/* out0069_em-eta9-phi3*/	7,37,0,9,37,1,9,37,2,5,93,1,2,93,2,3,94,1,3,94,2,4,
/* out0070_em-eta10-phi3*/	8,36,0,5,36,1,6,37,1,2,37,2,1,42,2,1,91,1,4,93,2,2,94,1,11,
/* out0071_em-eta11-phi3*/	5,36,0,11,36,2,1,41,1,2,91,1,5,91,2,8,
/* out0072_em-eta12-phi3*/	6,35,0,2,41,1,3,41,2,6,90,1,6,91,2,5,92,1,1,
/* out0073_em-eta13-phi3*/	6,35,0,3,40,1,4,41,2,3,90,0,3,90,1,5,90,2,2,
/* out0074_em-eta14-phi3*/	6,40,0,1,40,1,6,40,2,2,89,1,1,90,0,3,90,2,5,
/* out0075_em-eta15-phi3*/	4,40,2,6,89,0,4,89,1,2,96,2,1,
/* out0076_em-eta16-phi3*/	3,39,1,4,40,2,2,89,0,6,
/* out0077_em-eta17-phi3*/	3,39,1,4,89,0,2,95,1,4,
/* out0078_em-eta18-phi3*/	2,39,0,5,95,0,1,
/* out0079_em-eta19-phi3*/	0,
/* out0080_em-eta0-phi4*/	1,115,0,4,
/* out0081_em-eta1-phi4*/	2,114,0,6,115,0,12,
/* out0082_em-eta2-phi4*/	2,114,0,10,114,1,8,
/* out0083_em-eta3-phi4*/	2,113,0,9,114,1,8,
/* out0084_em-eta4-phi4*/	2,113,0,7,113,1,10,
/* out0085_em-eta5-phi4*/	2,112,0,11,113,1,6,
/* out0086_em-eta6-phi4*/	2,112,0,5,112,1,16,
/* out0087_em-eta7-phi4*/	0,
/* out0088_em-eta8-phi4*/	0,
/* out0089_em-eta9-phi4*/	6,37,0,1,37,1,5,38,0,7,38,2,11,94,0,1,94,2,11,
/* out0090_em-eta10-phi4*/	7,36,1,10,36,2,3,38,2,5,92,2,1,94,0,13,94,1,2,94,2,1,
/* out0091_em-eta11-phi4*/	5,35,1,1,36,2,12,92,1,6,92,2,7,94,0,1,
/* out0092_em-eta12-phi4*/	5,35,0,3,35,1,8,90,1,2,92,0,1,92,1,9,
/* out0093_em-eta13-phi4*/	5,35,0,7,35,2,2,90,1,2,90,2,5,100,1,2,
/* out0094_em-eta14-phi4*/	8,29,1,2,35,0,1,35,2,1,40,1,2,40,2,3,89,1,3,90,2,4,100,1,1,
/* out0095_em-eta15-phi4*/	3,29,1,3,40,2,3,89,1,7,
/* out0096_em-eta16-phi4*/	4,39,1,2,39,2,3,89,0,2,89,2,3,
/* out0097_em-eta17-phi4*/	5,39,0,2,39,1,2,39,2,3,89,0,1,89,2,3,
/* out0098_em-eta18-phi4*/	1,39,0,6,
/* out0099_em-eta19-phi4*/	0,
/* out0100_em-eta0-phi5*/	1,115,1,4,
/* out0101_em-eta1-phi5*/	2,114,3,6,115,1,12,
/* out0102_em-eta2-phi5*/	2,114,2,8,114,3,10,
/* out0103_em-eta3-phi5*/	2,113,3,9,114,2,8,
/* out0104_em-eta4-phi5*/	2,113,2,10,113,3,7,
/* out0105_em-eta5-phi5*/	2,112,3,11,113,2,6,
/* out0106_em-eta6-phi5*/	2,112,2,16,112,3,5,
/* out0107_em-eta7-phi5*/	0,
/* out0108_em-eta8-phi5*/	0,
/* out0109_em-eta9-phi5*/	4,38,0,9,38,1,10,102,0,1,102,1,6,
/* out0110_em-eta10-phi5*/	7,31,0,2,31,1,7,38,1,6,92,2,1,94,0,1,102,0,13,102,1,1,
/* out0111_em-eta11-phi5*/	5,31,0,13,35,1,1,92,0,5,92,2,7,102,0,2,
/* out0112_em-eta12-phi5*/	5,31,0,1,35,1,6,35,2,4,92,0,10,100,2,2,
/* out0113_em-eta13-phi5*/	4,29,2,1,35,2,9,100,1,4,100,2,6,
/* out0114_em-eta14-phi5*/	3,29,1,1,29,2,6,100,1,8,
/* out0115_em-eta15-phi5*/	4,29,1,7,89,1,3,89,2,2,100,1,1,
/* out0116_em-eta16-phi5*/	3,29,1,3,39,2,2,89,2,6,
/* out0117_em-eta17-phi5*/	2,39,2,5,89,2,2,
/* out0118_em-eta18-phi5*/	2,39,0,2,39,2,3,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	1,119,0,4,
/* out0121_em-eta1-phi6*/	2,118,0,6,119,0,12,
/* out0122_em-eta2-phi6*/	2,118,0,10,118,1,8,
/* out0123_em-eta3-phi6*/	2,117,0,9,118,1,8,
/* out0124_em-eta4-phi6*/	2,117,0,7,117,1,10,
/* out0125_em-eta5-phi6*/	2,116,0,11,117,1,6,
/* out0126_em-eta6-phi6*/	2,116,0,5,116,1,16,
/* out0127_em-eta7-phi6*/	0,
/* out0128_em-eta8-phi6*/	0,
/* out0129_em-eta9-phi6*/	5,33,0,11,33,1,2,33,2,10,102,1,7,102,2,1,
/* out0130_em-eta10-phi6*/	8,31,1,8,31,2,2,33,1,1,33,2,6,101,2,1,102,1,2,102,2,13,103,1,1,
/* out0131_em-eta11-phi6*/	6,30,2,1,31,1,1,31,2,13,101,1,5,101,2,7,102,2,2,
/* out0132_em-eta12-phi6*/	5,30,1,4,30,2,6,31,2,1,100,2,2,101,1,9,
/* out0133_em-eta13-phi6*/	4,29,2,1,30,1,9,100,0,4,100,2,6,
/* out0134_em-eta14-phi6*/	3,29,0,1,29,2,7,100,0,7,
/* out0135_em-eta15-phi6*/	4,29,0,6,85,1,2,85,2,3,100,0,1,
/* out0136_em-eta16-phi6*/	3,24,1,2,29,0,4,85,1,6,
/* out0137_em-eta17-phi6*/	2,24,1,4,85,1,2,
/* out0138_em-eta18-phi6*/	2,24,0,2,24,1,2,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	1,119,1,4,
/* out0141_em-eta1-phi7*/	2,118,3,6,119,1,12,
/* out0142_em-eta2-phi7*/	2,118,2,8,118,3,10,
/* out0143_em-eta3-phi7*/	2,117,3,9,118,2,8,
/* out0144_em-eta4-phi7*/	2,117,2,10,117,3,7,
/* out0145_em-eta5-phi7*/	2,116,3,11,117,2,6,
/* out0146_em-eta6-phi7*/	2,116,2,16,116,3,5,
/* out0147_em-eta7-phi7*/	0,
/* out0148_em-eta8-phi7*/	0,
/* out0149_em-eta9-phi7*/	6,33,0,5,33,1,10,34,0,2,34,2,5,103,1,1,103,2,11,
/* out0150_em-eta10-phi7*/	7,32,1,3,32,2,10,33,1,3,101,2,1,103,0,2,103,1,13,103,2,1,
/* out0151_em-eta11-phi7*/	5,30,2,1,32,1,12,101,0,6,101,2,7,103,1,1,
/* out0152_em-eta12-phi7*/	5,30,0,3,30,2,8,86,2,2,101,0,9,101,1,2,
/* out0153_em-eta13-phi7*/	5,30,0,7,30,1,2,86,1,5,86,2,2,100,0,2,
/* out0154_em-eta14-phi7*/	9,25,1,3,25,2,2,29,0,2,29,2,1,30,0,1,30,1,1,85,2,3,86,1,4,100,0,2,
/* out0155_em-eta15-phi7*/	3,25,1,3,29,0,3,85,2,7,
/* out0156_em-eta16-phi7*/	4,24,1,4,24,2,2,85,0,2,85,1,3,
/* out0157_em-eta17-phi7*/	4,24,0,1,24,1,4,85,0,1,85,1,3,
/* out0158_em-eta18-phi7*/	1,24,0,5,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	1,123,0,4,
/* out0161_em-eta1-phi8*/	2,122,0,6,123,0,12,
/* out0162_em-eta2-phi8*/	2,122,0,10,122,1,8,
/* out0163_em-eta3-phi8*/	2,121,0,9,122,1,8,
/* out0164_em-eta4-phi8*/	2,121,0,7,121,1,10,
/* out0165_em-eta5-phi8*/	2,120,0,11,121,1,6,
/* out0166_em-eta6-phi8*/	2,120,0,5,120,1,16,
/* out0167_em-eta7-phi8*/	0,
/* out0168_em-eta8-phi8*/	1,34,0,4,
/* out0169_em-eta9-phi8*/	7,34,0,9,34,1,7,34,2,8,88,1,3,88,2,2,103,0,3,103,2,4,
/* out0170_em-eta10-phi8*/	8,27,1,1,32,0,5,32,2,6,34,1,1,34,2,3,87,2,4,88,1,2,103,0,11,
/* out0171_em-eta11-phi8*/	5,26,2,2,32,0,11,32,1,1,87,1,8,87,2,5,
/* out0172_em-eta12-phi8*/	6,26,1,6,26,2,3,30,0,2,86,2,6,87,1,5,101,0,1,
/* out0173_em-eta13-phi8*/	6,25,2,4,26,1,3,30,0,3,86,0,3,86,1,2,86,2,5,
/* out0174_em-eta14-phi8*/	6,25,0,1,25,1,2,25,2,6,85,2,1,86,0,3,86,1,5,
/* out0175_em-eta15-phi8*/	4,25,1,6,81,1,1,85,0,4,85,2,2,
/* out0176_em-eta16-phi8*/	3,24,2,5,25,1,2,85,0,6,
/* out0177_em-eta17-phi8*/	4,24,0,2,24,2,4,80,1,4,85,0,2,
/* out0178_em-eta18-phi8*/	2,24,0,5,80,1,1,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	1,123,1,4,
/* out0181_em-eta1-phi9*/	2,122,3,6,123,1,12,
/* out0182_em-eta2-phi9*/	2,122,2,8,122,3,10,
/* out0183_em-eta3-phi9*/	2,121,3,9,122,2,8,
/* out0184_em-eta4-phi9*/	2,121,2,10,121,3,7,
/* out0185_em-eta5-phi9*/	2,120,3,11,121,2,6,
/* out0186_em-eta6-phi9*/	2,120,2,16,120,3,5,
/* out0187_em-eta7-phi9*/	0,
/* out0188_em-eta8-phi9*/	5,28,0,3,28,1,2,34,0,1,34,1,1,88,2,1,
/* out0189_em-eta9-phi9*/	6,27,2,5,28,1,10,34,1,7,88,0,5,88,1,3,88,2,13,
/* out0190_em-eta10-phi9*/	9,27,0,1,27,1,8,27,2,8,83,1,1,83,2,1,87,0,1,87,2,4,88,0,4,88,1,8,
/* out0191_em-eta11-phi9*/	5,26,2,7,27,1,6,87,0,11,87,1,1,87,2,3,
/* out0192_em-eta12-phi9*/	9,26,0,5,26,1,3,26,2,4,82,1,2,82,2,3,86,0,1,86,2,1,87,0,3,87,1,2,
/* out0193_em-eta13-phi9*/	5,25,2,2,26,0,2,26,1,4,82,1,3,86,0,6,
/* out0194_em-eta14-phi9*/	4,25,0,6,25,2,2,81,2,6,86,0,3,
/* out0195_em-eta15-phi9*/	3,25,0,6,81,1,5,81,2,2,
/* out0196_em-eta16-phi9*/	8,20,1,2,20,2,2,24,2,1,25,0,1,80,1,1,80,2,1,81,1,4,85,0,1,
/* out0197_em-eta17-phi9*/	4,20,1,2,24,2,3,80,1,4,80,2,2,
/* out0198_em-eta18-phi9*/	3,24,0,1,24,2,1,80,1,3,
/* out0199_em-eta19-phi9*/	0,
/* out0200_em-eta0-phi10*/	1,127,0,4,
/* out0201_em-eta1-phi10*/	2,126,0,6,127,0,12,
/* out0202_em-eta2-phi10*/	2,126,0,10,126,1,8,
/* out0203_em-eta3-phi10*/	2,125,0,9,126,1,8,
/* out0204_em-eta4-phi10*/	2,125,0,7,125,1,10,
/* out0205_em-eta5-phi10*/	2,124,0,11,125,1,6,
/* out0206_em-eta6-phi10*/	2,124,0,5,124,1,16,
/* out0207_em-eta7-phi10*/	0,
/* out0208_em-eta8-phi10*/	1,28,0,2,
/* out0209_em-eta9-phi10*/	9,23,1,2,23,2,4,27,0,1,27,2,2,28,0,11,28,1,4,84,0,3,84,1,13,88,0,5,
/* out0210_em-eta10-phi10*/	7,22,2,1,23,1,3,27,0,11,27,2,1,83,1,2,83,2,12,88,0,2,
/* out0211_em-eta11-phi10*/	8,22,1,3,22,2,5,26,0,1,27,0,3,27,1,1,82,2,2,83,1,11,87,0,1,
/* out0212_em-eta12-phi10*/	6,21,2,2,22,1,4,26,0,6,82,0,1,82,1,1,82,2,10,
/* out0213_em-eta13-phi10*/	5,21,1,1,21,2,7,26,0,2,82,0,1,82,1,9,
/* out0214_em-eta14-phi10*/	5,21,1,7,25,0,1,81,0,1,81,2,7,82,1,1,
/* out0215_em-eta15-phi10*/	6,20,2,5,21,1,1,25,0,1,81,0,3,81,1,2,81,2,1,
/* out0216_em-eta16-phi10*/	5,20,1,2,20,2,4,80,2,1,81,0,1,81,1,4,
/* out0217_em-eta17-phi10*/	2,20,1,5,80,2,7,
/* out0218_em-eta18-phi10*/	3,20,1,2,80,1,2,80,2,1,
/* out0219_em-eta19-phi10*/	0,
/* out0220_em-eta0-phi11*/	1,127,1,4,
/* out0221_em-eta1-phi11*/	2,126,3,6,127,1,12,
/* out0222_em-eta2-phi11*/	2,126,2,8,126,3,10,
/* out0223_em-eta3-phi11*/	2,125,3,9,126,2,8,
/* out0224_em-eta4-phi11*/	2,125,2,10,125,3,7,
/* out0225_em-eta5-phi11*/	2,124,3,11,125,2,6,
/* out0226_em-eta6-phi11*/	2,124,2,16,124,3,5,
/* out0227_em-eta7-phi11*/	0,
/* out0228_em-eta8-phi11*/	0,
/* out0229_em-eta9-phi11*/	6,23,0,5,23,1,2,23,2,12,79,0,3,84,0,13,84,1,3,
/* out0230_em-eta10-phi11*/	6,22,2,4,23,0,3,23,1,9,79,0,4,83,0,9,83,2,3,
/* out0231_em-eta11-phi11*/	6,22,0,6,22,1,2,22,2,6,78,0,4,83,0,7,83,1,2,
/* out0232_em-eta12-phi11*/	6,21,2,2,22,0,2,22,1,7,78,0,3,82,0,8,82,2,1,
/* out0233_em-eta13-phi11*/	4,21,0,5,21,2,5,77,0,3,82,0,6,
/* out0234_em-eta14-phi11*/	4,21,0,4,21,1,5,77,0,4,81,0,3,
/* out0235_em-eta15-phi11*/	4,20,0,1,20,2,4,21,1,2,81,0,6,
/* out0236_em-eta16-phi11*/	4,20,0,4,20,2,1,76,0,3,81,0,2,
/* out0237_em-eta17-phi11*/	4,20,0,3,20,1,2,76,0,3,80,2,2,
/* out0238_em-eta18-phi11*/	4,20,1,1,76,0,1,80,1,1,80,2,2,
/* out0239_em-eta19-phi11*/	0,
/* out0240_em-eta0-phi12*/	1,131,0,4,
/* out0241_em-eta1-phi12*/	2,130,0,6,131,0,12,
/* out0242_em-eta2-phi12*/	2,130,0,10,130,1,8,
/* out0243_em-eta3-phi12*/	2,129,0,9,130,1,8,
/* out0244_em-eta4-phi12*/	2,129,0,7,129,1,10,
/* out0245_em-eta5-phi12*/	2,128,0,11,129,1,6,
/* out0246_em-eta6-phi12*/	2,128,0,5,128,1,16,
/* out0247_em-eta7-phi12*/	0,
/* out0248_em-eta8-phi12*/	0,
/* out0249_em-eta9-phi12*/	6,18,1,1,19,0,13,19,2,4,23,0,5,79,0,4,79,1,12,
/* out0250_em-eta10-phi12*/	6,18,0,12,18,1,2,23,0,3,78,1,1,79,0,5,79,2,11,
/* out0251_em-eta11-phi12*/	7,17,0,1,17,1,1,18,0,4,18,2,2,22,0,6,78,0,5,78,1,9,
/* out0252_em-eta12-phi12*/	4,17,0,9,22,0,2,78,0,4,78,2,8,
/* out0253_em-eta13-phi12*/	5,17,0,4,17,2,1,21,0,4,77,0,3,77,1,7,
/* out0254_em-eta14-phi12*/	4,16,0,4,21,0,3,77,0,5,77,2,4,
/* out0255_em-eta15-phi12*/	6,16,0,6,20,0,1,76,0,1,76,1,3,77,0,1,77,2,3,
/* out0256_em-eta16-phi12*/	4,16,0,1,20,0,4,76,0,4,76,1,2,
/* out0257_em-eta17-phi12*/	4,15,0,3,20,0,3,76,0,3,76,2,1,
/* out0258_em-eta18-phi12*/	4,15,0,2,15,1,1,76,0,1,76,2,2,
/* out0259_em-eta19-phi12*/	0,
/* out0260_em-eta0-phi13*/	1,131,1,4,
/* out0261_em-eta1-phi13*/	2,130,3,6,131,1,12,
/* out0262_em-eta2-phi13*/	2,130,2,8,130,3,10,
/* out0263_em-eta3-phi13*/	2,129,3,9,130,2,8,
/* out0264_em-eta4-phi13*/	2,129,2,10,129,3,7,
/* out0265_em-eta5-phi13*/	2,128,3,11,129,2,6,
/* out0266_em-eta6-phi13*/	2,128,2,16,128,3,5,
/* out0267_em-eta7-phi13*/	0,
/* out0268_em-eta8-phi13*/	1,19,0,1,
/* out0269_em-eta9-phi13*/	8,14,0,7,18,1,3,19,0,2,19,2,12,74,1,1,75,0,13,75,2,4,79,1,4,
/* out0270_em-eta10-phi13*/	6,14,0,1,18,1,10,18,2,5,74,0,10,74,1,2,79,2,5,
/* out0271_em-eta11-phi13*/	8,12,0,1,17,1,5,18,2,8,73,0,1,74,0,5,74,2,1,78,1,6,78,2,2,
/* out0272_em-eta12-phi13*/	5,17,0,2,17,1,7,17,2,3,73,0,6,78,2,6,
/* out0273_em-eta13-phi13*/	4,16,1,1,17,2,8,73,0,2,77,1,8,
/* out0274_em-eta14-phi13*/	4,16,0,1,16,1,7,77,1,1,77,2,7,
/* out0275_em-eta15-phi13*/	6,16,0,3,16,1,1,16,2,3,72,0,1,76,1,4,77,2,2,
/* out0276_em-eta16-phi13*/	5,15,0,2,16,0,1,16,2,3,76,1,5,76,2,1,
/* out0277_em-eta17-phi13*/	2,15,0,6,76,2,5,
/* out0278_em-eta18-phi13*/	2,15,1,2,76,2,3,
/* out0279_em-eta19-phi13*/	0,
/* out0280_em-eta0-phi14*/	1,135,0,4,
/* out0281_em-eta1-phi14*/	2,134,0,6,135,0,12,
/* out0282_em-eta2-phi14*/	2,134,0,10,134,1,8,
/* out0283_em-eta3-phi14*/	2,133,0,9,134,1,8,
/* out0284_em-eta4-phi14*/	2,133,0,7,133,1,10,
/* out0285_em-eta5-phi14*/	2,132,0,11,133,1,6,
/* out0286_em-eta6-phi14*/	2,132,0,5,132,1,16,
/* out0287_em-eta7-phi14*/	0,
/* out0288_em-eta8-phi14*/	2,14,1,5,75,0,1,
/* out0289_em-eta9-phi14*/	8,14,0,6,14,1,9,14,2,5,70,0,1,70,2,9,74,1,2,75,0,2,75,2,12,
/* out0290_em-eta10-phi14*/	9,12,0,2,12,1,6,14,0,2,14,2,6,18,2,1,70,2,1,74,0,1,74,1,11,74,2,5,
/* out0291_em-eta11-phi14*/	5,12,0,11,12,1,1,12,2,1,73,1,5,74,2,9,
/* out0292_em-eta12-phi14*/	9,10,0,2,10,1,1,12,0,2,12,2,2,17,1,3,17,2,2,73,0,4,73,1,6,73,2,2,
/* out0293_em-eta13-phi14*/	6,10,0,7,16,1,1,17,2,2,72,1,1,73,0,3,73,2,6,
/* out0294_em-eta14-phi14*/	4,10,0,1,16,1,6,72,0,5,72,1,3,
/* out0295_em-eta15-phi14*/	2,16,2,6,72,0,7,
/* out0296_em-eta16-phi14*/	8,9,0,1,15,0,2,15,1,1,16,2,3,71,1,1,72,0,2,76,1,2,76,2,1,
/* out0297_em-eta17-phi14*/	4,15,0,1,15,1,5,71,1,2,76,2,2,
/* out0298_em-eta18-phi14*/	4,15,1,1,71,0,1,71,1,1,76,2,1,
/* out0299_em-eta19-phi14*/	0,
/* out0300_em-eta0-phi15*/	1,135,1,4,
/* out0301_em-eta1-phi15*/	2,134,3,6,135,1,12,
/* out0302_em-eta2-phi15*/	2,134,2,8,134,3,10,
/* out0303_em-eta3-phi15*/	2,133,3,9,134,2,8,
/* out0304_em-eta4-phi15*/	2,133,2,10,133,3,7,
/* out0305_em-eta5-phi15*/	2,132,3,11,133,2,6,
/* out0306_em-eta6-phi15*/	2,132,2,16,132,3,5,
/* out0307_em-eta7-phi15*/	0,
/* out0308_em-eta8-phi15*/	0,
/* out0309_em-eta9-phi15*/	7,13,1,5,13,2,4,14,1,2,14,2,4,70,0,14,70,1,7,70,2,4,
/* out0310_em-eta10-phi15*/	8,12,1,6,13,1,9,14,2,1,68,0,3,68,1,6,70,1,5,70,2,2,74,2,1,
/* out0311_em-eta11-phi15*/	5,11,1,1,12,1,3,12,2,10,68,0,12,73,1,1,
/* out0312_em-eta12-phi15*/	7,10,1,8,12,2,3,67,0,2,68,0,1,68,2,1,73,1,4,73,2,4,
/* out0313_em-eta13-phi15*/	6,10,0,4,10,1,3,10,2,3,67,0,3,72,1,2,73,2,4,
/* out0314_em-eta14-phi15*/	5,9,1,2,10,0,2,10,2,4,72,1,8,72,2,1,
/* out0315_em-eta15-phi15*/	5,9,0,5,9,1,1,16,2,1,72,0,1,72,2,6,
/* out0316_em-eta16-phi15*/	4,9,0,5,15,1,1,71,1,3,72,2,3,
/* out0317_em-eta17-phi15*/	3,9,0,1,15,1,5,71,1,4,
/* out0318_em-eta18-phi15*/	2,71,0,5,71,1,1,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	1,139,0,4,
/* out0321_em-eta1-phi16*/	2,138,0,6,139,0,12,
/* out0322_em-eta2-phi16*/	2,138,0,10,138,1,8,
/* out0323_em-eta3-phi16*/	2,137,0,9,138,1,8,
/* out0324_em-eta4-phi16*/	2,137,0,7,137,1,10,
/* out0325_em-eta5-phi16*/	2,136,0,11,137,1,6,
/* out0326_em-eta6-phi16*/	2,136,0,5,136,1,16,
/* out0327_em-eta7-phi16*/	0,
/* out0328_em-eta8-phi16*/	0,
/* out0329_em-eta9-phi16*/	6,13,0,3,13,2,12,69,0,7,69,2,8,70,0,1,70,1,3,
/* out0330_em-eta10-phi16*/	7,11,2,3,13,0,12,13,1,2,68,1,9,68,2,1,69,2,8,70,1,1,
/* out0331_em-eta11-phi16*/	4,11,1,8,11,2,5,68,1,1,68,2,13,
/* out0332_em-eta12-phi16*/	6,10,1,3,11,0,2,11,1,7,67,0,2,67,1,9,68,2,1,
/* out0333_em-eta13-phi16*/	6,10,1,1,10,2,6,48,1,2,67,0,7,67,1,1,67,2,2,
/* out0334_em-eta14-phi16*/	8,9,1,4,10,2,3,48,1,1,61,1,1,67,0,2,67,2,1,72,1,2,72,2,2,
/* out0335_em-eta15-phi16*/	5,9,0,1,9,1,5,9,2,1,61,1,3,72,2,4,
/* out0336_em-eta16-phi16*/	5,9,0,2,9,2,3,61,1,1,71,1,2,71,2,3,
/* out0337_em-eta17-phi16*/	4,9,0,1,9,2,2,71,1,2,71,2,3,
/* out0338_em-eta18-phi16*/	1,71,0,7,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	1,139,1,4,
/* out0341_em-eta1-phi17*/	2,138,3,6,139,1,12,
/* out0342_em-eta2-phi17*/	2,138,2,8,138,3,10,
/* out0343_em-eta3-phi17*/	2,137,3,9,138,2,8,
/* out0344_em-eta4-phi17*/	2,137,2,10,137,3,7,
/* out0345_em-eta5-phi17*/	2,136,3,11,137,2,6,
/* out0346_em-eta6-phi17*/	2,136,2,16,136,3,5,
/* out0347_em-eta7-phi17*/	0,
/* out0348_em-eta8-phi17*/	0,
/* out0349_em-eta9-phi17*/	5,13,0,1,51,0,3,51,1,8,69,0,9,69,1,7,
/* out0350_em-eta10-phi17*/	5,11,2,2,51,0,13,65,0,1,65,1,6,69,1,9,
/* out0351_em-eta11-phi17*/	4,11,0,7,11,2,6,65,0,12,65,1,2,
/* out0352_em-eta12-phi17*/	5,11,0,7,48,2,4,65,0,3,67,1,6,67,2,2,
/* out0353_em-eta13-phi17*/	3,48,1,6,48,2,4,67,2,10,
/* out0354_em-eta14-phi17*/	4,9,1,1,48,1,7,61,2,6,67,2,1,
/* out0355_em-eta15-phi17*/	4,9,1,3,9,2,4,61,1,6,61,2,1,
/* out0356_em-eta16-phi17*/	3,9,2,5,61,1,5,71,2,1,
/* out0357_em-eta17-phi17*/	2,9,2,1,71,2,6,
/* out0358_em-eta18-phi17*/	2,71,0,2,71,2,3,
/* out0359_em-eta19-phi17*/	1,71,0,1,
/* out0360_em-eta0-phi18*/	1,143,0,4,
/* out0361_em-eta1-phi18*/	2,142,0,6,143,0,12,
/* out0362_em-eta2-phi18*/	2,142,0,10,142,1,8,
/* out0363_em-eta3-phi18*/	2,141,0,9,142,1,8,
/* out0364_em-eta4-phi18*/	2,141,0,7,141,1,10,
/* out0365_em-eta5-phi18*/	2,140,0,11,141,1,6,
/* out0366_em-eta6-phi18*/	2,140,0,5,140,1,16,
/* out0367_em-eta7-phi18*/	0,
/* out0368_em-eta8-phi18*/	0,
/* out0369_em-eta9-phi18*/	6,50,1,1,51,1,8,51,2,3,66,0,11,66,1,1,66,2,7,
/* out0370_em-eta10-phi18*/	6,49,2,2,51,2,13,65,1,6,65,2,1,66,1,2,66,2,9,
/* out0371_em-eta11-phi18*/	4,49,1,7,49,2,6,65,1,2,65,2,12,
/* out0372_em-eta12-phi18*/	5,48,2,4,49,1,7,62,1,2,62,2,6,65,2,3,
/* out0373_em-eta13-phi18*/	3,48,0,6,48,2,4,62,1,10,
/* out0374_em-eta14-phi18*/	4,5,2,1,48,0,7,61,2,7,62,1,1,
/* out0375_em-eta15-phi18*/	4,5,1,4,5,2,3,61,0,6,61,2,1,
/* out0376_em-eta16-phi18*/	3,5,1,5,56,1,1,61,0,5,
/* out0377_em-eta17-phi18*/	2,5,1,1,56,1,4,
/* out0378_em-eta18-phi18*/	2,56,0,1,56,1,3,
/* out0379_em-eta19-phi18*/	1,56,0,1,
/* out0380_em-eta0-phi19*/	1,143,1,4,
/* out0381_em-eta1-phi19*/	2,142,3,6,143,1,12,
/* out0382_em-eta2-phi19*/	2,142,2,8,142,3,10,
/* out0383_em-eta3-phi19*/	2,141,3,9,142,2,8,
/* out0384_em-eta4-phi19*/	2,141,2,10,141,3,7,
/* out0385_em-eta5-phi19*/	2,140,3,11,141,2,6,
/* out0386_em-eta6-phi19*/	2,140,2,16,140,3,5,
/* out0387_em-eta7-phi19*/	0,
/* out0388_em-eta8-phi19*/	0,
/* out0389_em-eta9-phi19*/	6,50,1,3,50,2,12,64,0,2,64,2,5,66,0,5,66,1,7,
/* out0390_em-eta10-phi19*/	7,49,2,3,50,0,2,50,1,12,63,1,1,63,2,9,64,2,1,66,1,6,
/* out0391_em-eta11-phi19*/	4,49,0,8,49,2,5,63,1,13,63,2,1,
/* out0392_em-eta12-phi19*/	6,6,2,3,49,0,7,49,1,2,62,0,2,62,2,9,63,1,1,
/* out0393_em-eta13-phi19*/	6,6,1,6,6,2,1,48,0,2,62,0,7,62,1,2,62,2,1,
/* out0394_em-eta14-phi19*/	9,5,2,4,6,1,3,48,0,1,57,1,2,57,2,2,61,0,1,61,2,1,62,0,2,62,1,1,
/* out0395_em-eta15-phi19*/	5,5,0,1,5,1,1,5,2,5,57,1,4,61,0,3,
/* out0396_em-eta16-phi19*/	5,5,0,2,5,1,3,56,1,3,56,2,2,61,0,1,
/* out0397_em-eta17-phi19*/	3,5,0,1,5,1,2,56,1,4,
/* out0398_em-eta18-phi19*/	2,56,0,5,56,1,1,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	1,147,0,4,
/* out0401_em-eta1-phi20*/	2,146,0,6,147,0,12,
/* out0402_em-eta2-phi20*/	2,146,0,10,146,1,8,
/* out0403_em-eta3-phi20*/	2,145,0,9,146,1,8,
/* out0404_em-eta4-phi20*/	2,145,0,7,145,1,10,
/* out0405_em-eta5-phi20*/	2,144,0,11,145,1,6,
/* out0406_em-eta6-phi20*/	2,144,0,5,144,1,16,
/* out0407_em-eta7-phi20*/	0,
/* out0408_em-eta8-phi20*/	0,
/* out0409_em-eta9-phi20*/	7,8,1,4,8,2,2,50,0,5,50,2,4,64,0,14,64,1,6,64,2,5,
/* out0410_em-eta10-phi20*/	8,7,2,6,8,1,1,50,0,9,59,1,1,63,0,3,63,2,6,64,1,2,64,2,5,
/* out0411_em-eta11-phi20*/	5,7,1,10,7,2,3,49,0,1,58,2,1,63,0,12,
/* out0412_em-eta12-phi20*/	7,6,2,8,7,1,3,58,1,4,58,2,4,62,0,2,63,0,1,63,1,1,
/* out0413_em-eta13-phi20*/	6,6,0,4,6,1,3,6,2,3,57,2,2,58,1,4,62,0,3,
/* out0414_em-eta14-phi20*/	5,5,2,2,6,0,2,6,1,4,57,1,1,57,2,8,
/* out0415_em-eta15-phi20*/	5,1,1,1,5,0,5,5,2,1,57,0,1,57,1,6,
/* out0416_em-eta16-phi20*/	4,0,1,1,5,0,5,56,2,4,57,1,3,
/* out0417_em-eta17-phi20*/	4,0,1,5,5,0,1,56,0,1,56,2,5,
/* out0418_em-eta18-phi20*/	1,56,0,6,
/* out0419_em-eta19-phi20*/	0,
/* out0420_em-eta0-phi21*/	1,147,1,4,
/* out0421_em-eta1-phi21*/	2,146,3,6,147,1,12,
/* out0422_em-eta2-phi21*/	2,146,2,8,146,3,10,
/* out0423_em-eta3-phi21*/	2,145,3,9,146,2,8,
/* out0424_em-eta4-phi21*/	2,145,2,10,145,3,7,
/* out0425_em-eta5-phi21*/	2,144,3,11,145,2,6,
/* out0426_em-eta6-phi21*/	2,144,2,16,144,3,5,
/* out0427_em-eta7-phi21*/	0,
/* out0428_em-eta8-phi21*/	2,8,2,5,60,0,1,
/* out0429_em-eta9-phi21*/	7,8,0,6,8,1,5,8,2,9,59,2,2,60,0,2,60,1,12,64,1,7,
/* out0430_em-eta10-phi21*/	9,3,1,1,7,0,2,7,2,6,8,0,2,8,1,6,59,0,1,59,1,5,59,2,11,64,1,1,
/* out0431_em-eta11-phi21*/	5,7,0,11,7,1,1,7,2,1,58,2,5,59,1,9,
/* out0432_em-eta12-phi21*/	9,2,1,2,2,2,3,6,0,2,6,2,1,7,0,2,7,1,2,58,0,4,58,1,2,58,2,6,
/* out0433_em-eta13-phi21*/	6,1,2,1,2,1,2,6,0,7,57,2,1,58,0,3,58,1,6,
/* out0434_em-eta14-phi21*/	4,1,2,6,6,0,1,57,0,5,57,2,3,
/* out0435_em-eta15-phi21*/	2,1,1,6,57,0,7,
/* out0436_em-eta16-phi21*/	8,0,1,1,0,2,2,1,1,3,5,0,1,52,1,1,52,2,2,56,2,1,57,0,2,
/* out0437_em-eta17-phi21*/	4,0,1,5,0,2,1,52,1,2,56,2,3,
/* out0438_em-eta18-phi21*/	4,0,1,1,52,1,1,56,0,2,56,2,1,
/* out0439_em-eta19-phi21*/	0,
/* out0440_em-eta0-phi22*/	1,151,0,4,
/* out0441_em-eta1-phi22*/	2,150,0,6,151,0,12,
/* out0442_em-eta2-phi22*/	2,150,0,10,150,1,8,
/* out0443_em-eta3-phi22*/	2,149,0,9,150,1,8,
/* out0444_em-eta4-phi22*/	2,149,0,7,149,1,10,
/* out0445_em-eta5-phi22*/	2,148,0,11,149,1,6,
/* out0446_em-eta6-phi22*/	2,148,0,5,148,1,16,
/* out0447_em-eta7-phi22*/	0,
/* out0448_em-eta8-phi22*/	1,4,0,1,
/* out0449_em-eta9-phi22*/	8,3,2,3,4,0,2,4,1,12,8,0,7,55,2,4,59,2,1,60,0,13,60,1,4,
/* out0450_em-eta10-phi22*/	6,3,1,5,3,2,10,8,0,1,55,1,5,59,0,10,59,2,2,
/* out0451_em-eta11-phi22*/	8,2,2,5,3,1,8,7,0,1,54,1,2,54,2,6,58,0,1,59,0,5,59,1,1,
/* out0452_em-eta12-phi22*/	5,2,0,2,2,1,3,2,2,7,54,1,6,58,0,6,
/* out0453_em-eta13-phi22*/	4,1,2,1,2,1,8,53,2,8,58,0,2,
/* out0454_em-eta14-phi22*/	4,1,0,1,1,2,7,53,1,7,53,2,1,
/* out0455_em-eta15-phi22*/	6,1,0,3,1,1,3,1,2,1,52,2,4,53,1,2,57,0,1,
/* out0456_em-eta16-phi22*/	5,0,2,2,1,0,1,1,1,3,52,1,1,52,2,5,
/* out0457_em-eta17-phi22*/	2,0,2,6,52,1,5,
/* out0458_em-eta18-phi22*/	2,0,1,2,52,1,3,
/* out0459_em-eta19-phi22*/	0,
/* out0460_em-eta0-phi23*/	1,151,1,4,
/* out0461_em-eta1-phi23*/	2,150,3,6,151,1,12,
/* out0462_em-eta2-phi23*/	2,150,2,8,150,3,10,
/* out0463_em-eta3-phi23*/	2,149,3,9,150,2,8,
/* out0464_em-eta4-phi23*/	2,149,2,10,149,3,7,
/* out0465_em-eta5-phi23*/	2,148,3,11,149,2,6,
/* out0466_em-eta6-phi23*/	2,148,2,16,148,3,5,
/* out0467_em-eta7-phi23*/	0,
/* out0468_em-eta8-phi23*/	0,
/* out0469_em-eta9-phi23*/	5,3,2,1,4,0,13,4,1,4,55,0,4,55,2,12,
/* out0470_em-eta10-phi23*/	6,3,0,12,3,2,2,54,0,7,54,2,1,55,0,12,55,1,11,
/* out0471_em-eta11-phi23*/	6,2,0,1,2,2,1,3,0,4,3,1,2,54,0,5,54,2,9,
/* out0472_em-eta12-phi23*/	4,2,0,9,53,0,6,54,0,4,54,1,8,
/* out0473_em-eta13-phi23*/	4,2,0,4,2,1,1,53,0,4,53,2,7,
/* out0474_em-eta14-phi23*/	3,1,0,4,53,0,5,53,1,4,
/* out0475_em-eta15-phi23*/	5,1,0,6,52,0,1,52,2,3,53,0,1,53,1,3,
/* out0476_em-eta16-phi23*/	3,1,0,1,52,0,4,52,2,2,
/* out0477_em-eta17-phi23*/	3,0,2,3,52,0,10,52,1,1,
/* out0478_em-eta18-phi23*/	4,0,1,1,0,2,2,52,0,1,52,1,2,
/* out0479_em-eta19-phi23*/	0
};