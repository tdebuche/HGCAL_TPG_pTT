parameter integer matrixH [0:2612] = {
/* num inputs = 174(in0-in173) */
/* num outputs = 560(out0-out559) */
//* max inputs per outputs = 5 */
//* total number of input in adders 1026 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	1, 24, 1, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	1, 3, 1, 
/* out0033_had-eta13-phi1*/	1, 3, 1, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	1, 1, 1, 
/* out0036_had-eta16-phi1*/	1, 1, 1, 
/* out0037_had-eta17-phi1*/	1, 1, 1, 
/* out0038_had-eta18-phi1*/	1, 0, 1, 
/* out0039_had-eta19-phi1*/	1, 0, 2, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	1, 27, 2, 
/* out0045_had-eta5-phi2*/	1, 27, 5, 
/* out0046_had-eta6-phi2*/	1, 26, 6, 
/* out0047_had-eta7-phi2*/	2, 25, 2, 26, 2, 
/* out0048_had-eta8-phi2*/	1, 25, 5, 
/* out0049_had-eta9-phi2*/	2, 24, 2, 25, 1, 
/* out0050_had-eta10-phi2*/	1, 24, 4, 
/* out0051_had-eta11-phi2*/	2, 3, 1, 24, 1, 
/* out0052_had-eta12-phi2*/	1, 3, 2, 
/* out0053_had-eta13-phi2*/	1, 3, 2, 
/* out0054_had-eta14-phi2*/	2, 1, 1, 3, 1, 
/* out0055_had-eta15-phi2*/	1, 1, 2, 
/* out0056_had-eta16-phi2*/	1, 1, 1, 
/* out0057_had-eta17-phi2*/	1, 1, 1, 
/* out0058_had-eta18-phi2*/	1, 0, 2, 
/* out0059_had-eta19-phi2*/	1, 0, 2, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 118, 5, 
/* out0062_had-eta2-phi3*/	3, 36, 1, 117, 1, 118, 3, 
/* out0063_had-eta3-phi3*/	2, 36, 6, 117, 5, 
/* out0064_had-eta4-phi3*/	4, 27, 3, 35, 5, 116, 2, 117, 2, 
/* out0065_had-eta5-phi3*/	3, 27, 6, 34, 3, 116, 4, 
/* out0066_had-eta6-phi3*/	5, 26, 6, 33, 1, 34, 1, 115, 2, 116, 2, 
/* out0067_had-eta7-phi3*/	4, 25, 2, 26, 2, 33, 2, 115, 3, 
/* out0068_had-eta8-phi3*/	2, 25, 5, 115, 2, 
/* out0069_had-eta9-phi3*/	5, 24, 2, 25, 1, 32, 1, 114, 3, 115, 1, 
/* out0070_had-eta10-phi3*/	2, 24, 4, 114, 5, 
/* out0071_had-eta11-phi3*/	2, 3, 1, 24, 1, 
/* out0072_had-eta12-phi3*/	1, 3, 2, 
/* out0073_had-eta13-phi3*/	1, 3, 2, 
/* out0074_had-eta14-phi3*/	2, 1, 1, 3, 1, 
/* out0075_had-eta15-phi3*/	1, 1, 2, 
/* out0076_had-eta16-phi3*/	1, 1, 1, 
/* out0077_had-eta17-phi3*/	1, 1, 1, 
/* out0078_had-eta18-phi3*/	1, 0, 2, 
/* out0079_had-eta19-phi3*/	1, 0, 2, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 118, 5, 
/* out0082_had-eta2-phi4*/	3, 36, 1, 117, 1, 118, 3, 
/* out0083_had-eta3-phi4*/	4, 35, 1, 36, 8, 46, 4, 117, 5, 
/* out0084_had-eta4-phi4*/	5, 35, 9, 45, 1, 46, 1, 116, 2, 117, 2, 
/* out0085_had-eta5-phi4*/	4, 34, 7, 35, 1, 45, 1, 116, 4, 
/* out0086_had-eta6-phi4*/	4, 33, 3, 34, 4, 115, 2, 116, 2, 
/* out0087_had-eta7-phi4*/	2, 33, 6, 115, 3, 
/* out0088_had-eta8-phi4*/	3, 32, 4, 33, 1, 115, 2, 
/* out0089_had-eta9-phi4*/	3, 32, 4, 114, 3, 115, 1, 
/* out0090_had-eta10-phi4*/	4, 5, 2, 24, 1, 32, 1, 114, 5, 
/* out0091_had-eta11-phi4*/	1, 5, 3, 
/* out0092_had-eta12-phi4*/	2, 3, 1, 5, 1, 
/* out0093_had-eta13-phi4*/	2, 3, 1, 4, 1, 
/* out0094_had-eta14-phi4*/	1, 4, 1, 
/* out0095_had-eta15-phi4*/	1, 1, 1, 
/* out0096_had-eta16-phi4*/	1, 1, 1, 
/* out0097_had-eta17-phi4*/	1, 1, 1, 
/* out0098_had-eta18-phi4*/	1, 0, 2, 
/* out0099_had-eta19-phi4*/	1, 0, 2, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 123, 5, 
/* out0102_had-eta2-phi5*/	2, 122, 1, 123, 3, 
/* out0103_had-eta3-phi5*/	4, 46, 8, 55, 1, 56, 6, 122, 5, 
/* out0104_had-eta4-phi5*/	5, 45, 7, 46, 3, 55, 1, 121, 2, 122, 2, 
/* out0105_had-eta5-phi5*/	4, 34, 1, 44, 3, 45, 6, 121, 4, 
/* out0106_had-eta6-phi5*/	4, 33, 1, 44, 7, 120, 2, 121, 2, 
/* out0107_had-eta7-phi5*/	4, 33, 2, 43, 3, 44, 1, 120, 3, 
/* out0108_had-eta8-phi5*/	3, 32, 3, 43, 3, 120, 2, 
/* out0109_had-eta9-phi5*/	4, 32, 3, 42, 1, 119, 3, 120, 1, 
/* out0110_had-eta10-phi5*/	2, 5, 3, 119, 5, 
/* out0111_had-eta11-phi5*/	1, 5, 3, 
/* out0112_had-eta12-phi5*/	2, 4, 1, 5, 2, 
/* out0113_had-eta13-phi5*/	1, 4, 2, 
/* out0114_had-eta14-phi5*/	1, 4, 2, 
/* out0115_had-eta15-phi5*/	1, 4, 1, 
/* out0116_had-eta16-phi5*/	1, 2, 1, 
/* out0117_had-eta17-phi5*/	1, 2, 1, 
/* out0118_had-eta18-phi5*/	1, 2, 1, 
/* out0119_had-eta19-phi5*/	1, 0, 1, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 123, 5, 
/* out0122_had-eta2-phi6*/	4, 56, 1, 108, 1, 122, 1, 123, 3, 
/* out0123_had-eta3-phi6*/	4, 55, 6, 56, 9, 108, 4, 122, 5, 
/* out0124_had-eta4-phi6*/	5, 45, 1, 54, 3, 55, 8, 121, 2, 122, 2, 
/* out0125_had-eta5-phi6*/	3, 44, 1, 54, 8, 121, 4, 
/* out0126_had-eta6-phi6*/	4, 44, 4, 53, 3, 120, 2, 121, 2, 
/* out0127_had-eta7-phi6*/	3, 43, 5, 53, 1, 120, 3, 
/* out0128_had-eta8-phi6*/	3, 42, 1, 43, 4, 120, 2, 
/* out0129_had-eta9-phi6*/	3, 42, 4, 119, 3, 120, 1, 
/* out0130_had-eta10-phi6*/	3, 5, 1, 42, 3, 119, 5, 
/* out0131_had-eta11-phi6*/	2, 5, 1, 6, 2, 
/* out0132_had-eta12-phi6*/	2, 4, 1, 6, 1, 
/* out0133_had-eta13-phi6*/	1, 4, 2, 
/* out0134_had-eta14-phi6*/	1, 4, 2, 
/* out0135_had-eta15-phi6*/	2, 2, 1, 4, 1, 
/* out0136_had-eta16-phi6*/	1, 2, 1, 
/* out0137_had-eta17-phi6*/	1, 2, 1, 
/* out0138_had-eta18-phi6*/	1, 2, 1, 
/* out0139_had-eta19-phi6*/	1, 2, 1, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 128, 5, 
/* out0142_had-eta2-phi7*/	3, 108, 1, 127, 1, 128, 3, 
/* out0143_had-eta3-phi7*/	4, 107, 3, 108, 10, 109, 2, 127, 5, 
/* out0144_had-eta4-phi7*/	4, 54, 1, 107, 10, 126, 2, 127, 2, 
/* out0145_had-eta5-phi7*/	4, 53, 1, 54, 4, 106, 4, 126, 4, 
/* out0146_had-eta6-phi7*/	3, 53, 7, 125, 2, 126, 2, 
/* out0147_had-eta7-phi7*/	4, 43, 1, 52, 3, 53, 3, 125, 3, 
/* out0148_had-eta8-phi7*/	3, 42, 1, 52, 5, 125, 2, 
/* out0149_had-eta9-phi7*/	3, 42, 4, 124, 3, 125, 1, 
/* out0150_had-eta10-phi7*/	3, 6, 1, 42, 2, 124, 5, 
/* out0151_had-eta11-phi7*/	1, 6, 3, 
/* out0152_had-eta12-phi7*/	1, 6, 3, 
/* out0153_had-eta13-phi7*/	3, 4, 1, 6, 1, 7, 1, 
/* out0154_had-eta14-phi7*/	2, 4, 1, 7, 1, 
/* out0155_had-eta15-phi7*/	2, 2, 1, 7, 1, 
/* out0156_had-eta16-phi7*/	1, 2, 1, 
/* out0157_had-eta17-phi7*/	1, 2, 1, 
/* out0158_had-eta18-phi7*/	1, 2, 1, 
/* out0159_had-eta19-phi7*/	1, 2, 1, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 128, 5, 
/* out0162_had-eta2-phi8*/	3, 109, 2, 127, 1, 128, 3, 
/* out0163_had-eta3-phi8*/	3, 96, 1, 109, 12, 127, 5, 
/* out0164_had-eta4-phi8*/	5, 96, 7, 106, 2, 107, 3, 126, 2, 127, 2, 
/* out0165_had-eta5-phi8*/	2, 106, 9, 126, 4, 
/* out0166_had-eta6-phi8*/	5, 53, 1, 94, 5, 106, 1, 125, 2, 126, 2, 
/* out0167_had-eta7-phi8*/	3, 52, 3, 94, 3, 125, 3, 
/* out0168_had-eta8-phi8*/	2, 52, 5, 125, 2, 
/* out0169_had-eta9-phi8*/	3, 62, 4, 124, 3, 125, 1, 
/* out0170_had-eta10-phi8*/	2, 62, 3, 124, 5, 
/* out0171_had-eta11-phi8*/	1, 6, 3, 
/* out0172_had-eta12-phi8*/	1, 6, 2, 
/* out0173_had-eta13-phi8*/	1, 7, 2, 
/* out0174_had-eta14-phi8*/	1, 7, 2, 
/* out0175_had-eta15-phi8*/	1, 7, 1, 
/* out0176_had-eta16-phi8*/	1, 2, 1, 
/* out0177_had-eta17-phi8*/	1, 2, 1, 
/* out0178_had-eta18-phi8*/	1, 2, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 133, 5, 
/* out0182_had-eta2-phi9*/	3, 98, 2, 132, 1, 133, 3, 
/* out0183_had-eta3-phi9*/	3, 96, 1, 98, 12, 132, 5, 
/* out0184_had-eta4-phi9*/	5, 95, 2, 96, 7, 97, 3, 131, 2, 132, 2, 
/* out0185_had-eta5-phi9*/	2, 95, 9, 131, 4, 
/* out0186_had-eta6-phi9*/	5, 64, 1, 94, 5, 95, 1, 130, 2, 131, 2, 
/* out0187_had-eta7-phi9*/	3, 63, 3, 94, 3, 130, 3, 
/* out0188_had-eta8-phi9*/	2, 63, 5, 130, 2, 
/* out0189_had-eta9-phi9*/	3, 62, 4, 129, 3, 130, 1, 
/* out0190_had-eta10-phi9*/	2, 62, 3, 129, 5, 
/* out0191_had-eta11-phi9*/	1, 8, 3, 
/* out0192_had-eta12-phi9*/	1, 8, 2, 
/* out0193_had-eta13-phi9*/	1, 7, 2, 
/* out0194_had-eta14-phi9*/	1, 7, 2, 
/* out0195_had-eta15-phi9*/	1, 7, 1, 
/* out0196_had-eta16-phi9*/	1, 9, 1, 
/* out0197_had-eta17-phi9*/	1, 9, 1, 
/* out0198_had-eta18-phi9*/	1, 9, 1, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 133, 5, 
/* out0202_had-eta2-phi10*/	3, 99, 1, 132, 1, 133, 3, 
/* out0203_had-eta3-phi10*/	4, 97, 3, 98, 2, 99, 10, 132, 5, 
/* out0204_had-eta4-phi10*/	4, 65, 1, 97, 10, 131, 2, 132, 2, 
/* out0205_had-eta5-phi10*/	4, 64, 1, 65, 4, 95, 4, 131, 4, 
/* out0206_had-eta6-phi10*/	3, 64, 7, 130, 2, 131, 2, 
/* out0207_had-eta7-phi10*/	4, 63, 3, 64, 3, 75, 1, 130, 3, 
/* out0208_had-eta8-phi10*/	3, 63, 5, 74, 1, 130, 2, 
/* out0209_had-eta9-phi10*/	4, 62, 1, 74, 4, 129, 3, 130, 1, 
/* out0210_had-eta10-phi10*/	4, 8, 1, 62, 1, 74, 2, 129, 5, 
/* out0211_had-eta11-phi10*/	1, 8, 3, 
/* out0212_had-eta12-phi10*/	1, 8, 3, 
/* out0213_had-eta13-phi10*/	3, 7, 1, 8, 1, 10, 1, 
/* out0214_had-eta14-phi10*/	2, 7, 1, 10, 1, 
/* out0215_had-eta15-phi10*/	2, 7, 1, 9, 1, 
/* out0216_had-eta16-phi10*/	1, 9, 1, 
/* out0217_had-eta17-phi10*/	1, 9, 1, 
/* out0218_had-eta18-phi10*/	1, 9, 1, 
/* out0219_had-eta19-phi10*/	1, 9, 1, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 138, 5, 
/* out0222_had-eta2-phi11*/	4, 67, 1, 99, 1, 137, 1, 138, 3, 
/* out0223_had-eta3-phi11*/	4, 66, 6, 67, 9, 99, 4, 137, 5, 
/* out0224_had-eta4-phi11*/	5, 65, 3, 66, 8, 77, 1, 136, 2, 137, 2, 
/* out0225_had-eta5-phi11*/	3, 65, 8, 76, 1, 136, 4, 
/* out0226_had-eta6-phi11*/	4, 64, 3, 76, 4, 135, 2, 136, 2, 
/* out0227_had-eta7-phi11*/	3, 64, 1, 75, 5, 135, 3, 
/* out0228_had-eta8-phi11*/	3, 74, 1, 75, 4, 135, 2, 
/* out0229_had-eta9-phi11*/	3, 74, 4, 134, 3, 135, 1, 
/* out0230_had-eta10-phi11*/	3, 11, 1, 74, 3, 134, 5, 
/* out0231_had-eta11-phi11*/	2, 8, 2, 11, 1, 
/* out0232_had-eta12-phi11*/	2, 8, 1, 10, 1, 
/* out0233_had-eta13-phi11*/	1, 10, 2, 
/* out0234_had-eta14-phi11*/	1, 10, 2, 
/* out0235_had-eta15-phi11*/	2, 9, 1, 10, 1, 
/* out0236_had-eta16-phi11*/	1, 9, 1, 
/* out0237_had-eta17-phi11*/	1, 9, 1, 
/* out0238_had-eta18-phi11*/	1, 9, 1, 
/* out0239_had-eta19-phi11*/	1, 9, 1, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 138, 5, 
/* out0242_had-eta2-phi12*/	2, 137, 1, 138, 3, 
/* out0243_had-eta3-phi12*/	4, 66, 1, 67, 6, 78, 8, 137, 5, 
/* out0244_had-eta4-phi12*/	5, 66, 1, 77, 7, 78, 3, 136, 2, 137, 2, 
/* out0245_had-eta5-phi12*/	4, 76, 3, 77, 6, 86, 1, 136, 4, 
/* out0246_had-eta6-phi12*/	4, 76, 7, 85, 1, 135, 2, 136, 2, 
/* out0247_had-eta7-phi12*/	4, 75, 3, 76, 1, 85, 2, 135, 3, 
/* out0248_had-eta8-phi12*/	3, 75, 3, 84, 3, 135, 2, 
/* out0249_had-eta9-phi12*/	4, 74, 1, 84, 3, 134, 3, 135, 1, 
/* out0250_had-eta10-phi12*/	2, 11, 3, 134, 5, 
/* out0251_had-eta11-phi12*/	1, 11, 3, 
/* out0252_had-eta12-phi12*/	2, 10, 1, 11, 2, 
/* out0253_had-eta13-phi12*/	1, 10, 2, 
/* out0254_had-eta14-phi12*/	1, 10, 2, 
/* out0255_had-eta15-phi12*/	1, 10, 1, 
/* out0256_had-eta16-phi12*/	1, 9, 1, 
/* out0257_had-eta17-phi12*/	1, 9, 1, 
/* out0258_had-eta18-phi12*/	1, 9, 1, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 143, 5, 
/* out0262_had-eta2-phi13*/	3, 88, 1, 142, 1, 143, 3, 
/* out0263_had-eta3-phi13*/	4, 78, 4, 87, 1, 88, 8, 142, 5, 
/* out0264_had-eta4-phi13*/	5, 77, 1, 78, 1, 87, 9, 141, 2, 142, 2, 
/* out0265_had-eta5-phi13*/	4, 77, 1, 86, 7, 87, 1, 141, 4, 
/* out0266_had-eta6-phi13*/	4, 85, 3, 86, 4, 140, 2, 141, 2, 
/* out0267_had-eta7-phi13*/	2, 85, 6, 140, 3, 
/* out0268_had-eta8-phi13*/	3, 84, 4, 85, 1, 140, 2, 
/* out0269_had-eta9-phi13*/	3, 84, 4, 139, 3, 140, 1, 
/* out0270_had-eta10-phi13*/	4, 11, 2, 28, 1, 84, 1, 139, 5, 
/* out0271_had-eta11-phi13*/	1, 11, 3, 
/* out0272_had-eta12-phi13*/	2, 11, 1, 15, 1, 
/* out0273_had-eta13-phi13*/	2, 10, 1, 15, 1, 
/* out0274_had-eta14-phi13*/	1, 10, 1, 
/* out0275_had-eta15-phi13*/	1, 14, 1, 
/* out0276_had-eta16-phi13*/	1, 14, 1, 
/* out0277_had-eta17-phi13*/	1, 14, 1, 
/* out0278_had-eta18-phi13*/	1, 12, 1, 
/* out0279_had-eta19-phi13*/	1, 12, 2, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 143, 5, 
/* out0282_had-eta2-phi14*/	3, 88, 1, 142, 1, 143, 3, 
/* out0283_had-eta3-phi14*/	2, 88, 6, 142, 5, 
/* out0284_had-eta4-phi14*/	4, 31, 2, 87, 5, 141, 2, 142, 2, 
/* out0285_had-eta5-phi14*/	3, 31, 5, 86, 3, 141, 4, 
/* out0286_had-eta6-phi14*/	5, 30, 6, 85, 1, 86, 1, 140, 2, 141, 2, 
/* out0287_had-eta7-phi14*/	4, 29, 2, 30, 2, 85, 2, 140, 3, 
/* out0288_had-eta8-phi14*/	2, 29, 5, 140, 2, 
/* out0289_had-eta9-phi14*/	5, 28, 2, 29, 1, 84, 1, 139, 3, 140, 1, 
/* out0290_had-eta10-phi14*/	2, 28, 4, 139, 5, 
/* out0291_had-eta11-phi14*/	2, 15, 1, 28, 1, 
/* out0292_had-eta12-phi14*/	1, 15, 2, 
/* out0293_had-eta13-phi14*/	1, 15, 2, 
/* out0294_had-eta14-phi14*/	2, 14, 1, 15, 1, 
/* out0295_had-eta15-phi14*/	1, 14, 2, 
/* out0296_had-eta16-phi14*/	1, 14, 1, 
/* out0297_had-eta17-phi14*/	1, 14, 1, 
/* out0298_had-eta18-phi14*/	1, 12, 2, 
/* out0299_had-eta19-phi14*/	1, 12, 2, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 148, 5, 
/* out0302_had-eta2-phi15*/	3, 41, 1, 147, 1, 148, 3, 
/* out0303_had-eta3-phi15*/	2, 41, 6, 147, 5, 
/* out0304_had-eta4-phi15*/	4, 31, 3, 40, 5, 146, 2, 147, 2, 
/* out0305_had-eta5-phi15*/	3, 31, 6, 39, 3, 146, 4, 
/* out0306_had-eta6-phi15*/	5, 30, 6, 38, 1, 39, 1, 145, 2, 146, 2, 
/* out0307_had-eta7-phi15*/	4, 29, 2, 30, 2, 38, 2, 145, 3, 
/* out0308_had-eta8-phi15*/	2, 29, 5, 145, 2, 
/* out0309_had-eta9-phi15*/	5, 28, 2, 29, 1, 37, 1, 144, 3, 145, 1, 
/* out0310_had-eta10-phi15*/	2, 28, 4, 144, 5, 
/* out0311_had-eta11-phi15*/	2, 15, 1, 28, 1, 
/* out0312_had-eta12-phi15*/	1, 15, 2, 
/* out0313_had-eta13-phi15*/	1, 15, 2, 
/* out0314_had-eta14-phi15*/	2, 14, 1, 15, 1, 
/* out0315_had-eta15-phi15*/	1, 14, 2, 
/* out0316_had-eta16-phi15*/	1, 14, 1, 
/* out0317_had-eta17-phi15*/	1, 14, 1, 
/* out0318_had-eta18-phi15*/	1, 12, 2, 
/* out0319_had-eta19-phi15*/	1, 12, 2, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 148, 5, 
/* out0322_had-eta2-phi16*/	3, 41, 1, 147, 1, 148, 3, 
/* out0323_had-eta3-phi16*/	4, 40, 1, 41, 8, 51, 4, 147, 5, 
/* out0324_had-eta4-phi16*/	5, 40, 9, 50, 1, 51, 1, 146, 2, 147, 2, 
/* out0325_had-eta5-phi16*/	4, 39, 7, 40, 1, 50, 1, 146, 4, 
/* out0326_had-eta6-phi16*/	4, 38, 3, 39, 4, 145, 2, 146, 2, 
/* out0327_had-eta7-phi16*/	2, 38, 6, 145, 3, 
/* out0328_had-eta8-phi16*/	3, 37, 4, 38, 1, 145, 2, 
/* out0329_had-eta9-phi16*/	3, 37, 4, 144, 3, 145, 1, 
/* out0330_had-eta10-phi16*/	4, 18, 2, 28, 1, 37, 1, 144, 5, 
/* out0331_had-eta11-phi16*/	1, 18, 3, 
/* out0332_had-eta12-phi16*/	2, 15, 1, 18, 1, 
/* out0333_had-eta13-phi16*/	2, 15, 1, 16, 1, 
/* out0334_had-eta14-phi16*/	1, 16, 1, 
/* out0335_had-eta15-phi16*/	1, 14, 1, 
/* out0336_had-eta16-phi16*/	1, 14, 1, 
/* out0337_had-eta17-phi16*/	1, 14, 1, 
/* out0338_had-eta18-phi16*/	1, 12, 2, 
/* out0339_had-eta19-phi16*/	1, 12, 2, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 153, 5, 
/* out0342_had-eta2-phi17*/	2, 152, 1, 153, 3, 
/* out0343_had-eta3-phi17*/	4, 51, 8, 60, 1, 61, 6, 152, 5, 
/* out0344_had-eta4-phi17*/	5, 50, 7, 51, 3, 60, 1, 151, 2, 152, 2, 
/* out0345_had-eta5-phi17*/	4, 39, 1, 49, 3, 50, 6, 151, 4, 
/* out0346_had-eta6-phi17*/	4, 38, 1, 49, 7, 150, 2, 151, 2, 
/* out0347_had-eta7-phi17*/	4, 38, 2, 48, 3, 49, 1, 150, 3, 
/* out0348_had-eta8-phi17*/	3, 37, 3, 48, 3, 150, 2, 
/* out0349_had-eta9-phi17*/	4, 37, 3, 47, 1, 149, 3, 150, 1, 
/* out0350_had-eta10-phi17*/	2, 18, 3, 149, 5, 
/* out0351_had-eta11-phi17*/	1, 18, 3, 
/* out0352_had-eta12-phi17*/	2, 16, 1, 18, 2, 
/* out0353_had-eta13-phi17*/	1, 16, 2, 
/* out0354_had-eta14-phi17*/	1, 16, 2, 
/* out0355_had-eta15-phi17*/	1, 16, 1, 
/* out0356_had-eta16-phi17*/	1, 13, 1, 
/* out0357_had-eta17-phi17*/	1, 13, 1, 
/* out0358_had-eta18-phi17*/	1, 13, 1, 
/* out0359_had-eta19-phi17*/	1, 12, 1, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 153, 5, 
/* out0362_had-eta2-phi18*/	4, 61, 1, 113, 1, 152, 1, 153, 3, 
/* out0363_had-eta3-phi18*/	4, 60, 6, 61, 9, 113, 4, 152, 5, 
/* out0364_had-eta4-phi18*/	5, 50, 1, 59, 3, 60, 8, 151, 2, 152, 2, 
/* out0365_had-eta5-phi18*/	3, 49, 1, 59, 8, 151, 4, 
/* out0366_had-eta6-phi18*/	4, 49, 4, 58, 3, 150, 2, 151, 2, 
/* out0367_had-eta7-phi18*/	3, 48, 5, 58, 1, 150, 3, 
/* out0368_had-eta8-phi18*/	3, 47, 1, 48, 4, 150, 2, 
/* out0369_had-eta9-phi18*/	3, 47, 4, 149, 3, 150, 1, 
/* out0370_had-eta10-phi18*/	3, 18, 1, 47, 3, 149, 5, 
/* out0371_had-eta11-phi18*/	2, 17, 2, 18, 1, 
/* out0372_had-eta12-phi18*/	2, 16, 1, 17, 1, 
/* out0373_had-eta13-phi18*/	1, 16, 2, 
/* out0374_had-eta14-phi18*/	1, 16, 2, 
/* out0375_had-eta15-phi18*/	2, 13, 1, 16, 1, 
/* out0376_had-eta16-phi18*/	1, 13, 1, 
/* out0377_had-eta17-phi18*/	1, 13, 1, 
/* out0378_had-eta18-phi18*/	1, 13, 1, 
/* out0379_had-eta19-phi18*/	1, 13, 1, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 158, 5, 
/* out0382_had-eta2-phi19*/	3, 113, 1, 157, 1, 158, 3, 
/* out0383_had-eta3-phi19*/	4, 111, 3, 112, 2, 113, 10, 157, 5, 
/* out0384_had-eta4-phi19*/	4, 59, 1, 111, 10, 156, 2, 157, 2, 
/* out0385_had-eta5-phi19*/	4, 58, 1, 59, 4, 110, 4, 156, 4, 
/* out0386_had-eta6-phi19*/	3, 58, 7, 155, 2, 156, 2, 
/* out0387_had-eta7-phi19*/	4, 48, 1, 57, 3, 58, 3, 155, 3, 
/* out0388_had-eta8-phi19*/	3, 47, 1, 57, 5, 155, 2, 
/* out0389_had-eta9-phi19*/	3, 47, 4, 154, 3, 155, 1, 
/* out0390_had-eta10-phi19*/	3, 17, 1, 47, 2, 154, 5, 
/* out0391_had-eta11-phi19*/	1, 17, 3, 
/* out0392_had-eta12-phi19*/	1, 17, 3, 
/* out0393_had-eta13-phi19*/	3, 16, 1, 17, 1, 19, 1, 
/* out0394_had-eta14-phi19*/	2, 16, 1, 19, 1, 
/* out0395_had-eta15-phi19*/	2, 13, 1, 19, 1, 
/* out0396_had-eta16-phi19*/	1, 13, 1, 
/* out0397_had-eta17-phi19*/	1, 13, 1, 
/* out0398_had-eta18-phi19*/	1, 13, 1, 
/* out0399_had-eta19-phi19*/	1, 13, 1, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 158, 5, 
/* out0402_had-eta2-phi20*/	3, 112, 2, 157, 1, 158, 3, 
/* out0403_had-eta3-phi20*/	3, 104, 1, 112, 12, 157, 5, 
/* out0404_had-eta4-phi20*/	5, 104, 7, 110, 2, 111, 3, 156, 2, 157, 2, 
/* out0405_had-eta5-phi20*/	2, 110, 9, 156, 4, 
/* out0406_had-eta6-phi20*/	5, 58, 1, 100, 5, 110, 1, 155, 2, 156, 2, 
/* out0407_had-eta7-phi20*/	3, 57, 3, 100, 3, 155, 3, 
/* out0408_had-eta8-phi20*/	2, 57, 5, 155, 2, 
/* out0409_had-eta9-phi20*/	3, 68, 4, 154, 3, 155, 1, 
/* out0410_had-eta10-phi20*/	2, 68, 3, 154, 5, 
/* out0411_had-eta11-phi20*/	1, 17, 3, 
/* out0412_had-eta12-phi20*/	1, 17, 2, 
/* out0413_had-eta13-phi20*/	1, 19, 2, 
/* out0414_had-eta14-phi20*/	1, 19, 2, 
/* out0415_had-eta15-phi20*/	1, 19, 1, 
/* out0416_had-eta16-phi20*/	1, 13, 1, 
/* out0417_had-eta17-phi20*/	1, 13, 1, 
/* out0418_had-eta18-phi20*/	1, 13, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 163, 5, 
/* out0422_had-eta2-phi21*/	3, 105, 2, 162, 1, 163, 3, 
/* out0423_had-eta3-phi21*/	3, 104, 1, 105, 12, 162, 5, 
/* out0424_had-eta4-phi21*/	5, 101, 2, 102, 3, 104, 7, 161, 2, 162, 2, 
/* out0425_had-eta5-phi21*/	2, 101, 9, 161, 4, 
/* out0426_had-eta6-phi21*/	5, 70, 1, 100, 5, 101, 1, 160, 2, 161, 2, 
/* out0427_had-eta7-phi21*/	3, 69, 3, 100, 3, 160, 3, 
/* out0428_had-eta8-phi21*/	2, 69, 5, 160, 2, 
/* out0429_had-eta9-phi21*/	3, 68, 4, 159, 3, 160, 1, 
/* out0430_had-eta10-phi21*/	2, 68, 3, 159, 5, 
/* out0431_had-eta11-phi21*/	1, 20, 3, 
/* out0432_had-eta12-phi21*/	1, 20, 2, 
/* out0433_had-eta13-phi21*/	1, 19, 2, 
/* out0434_had-eta14-phi21*/	1, 19, 2, 
/* out0435_had-eta15-phi21*/	1, 19, 1, 
/* out0436_had-eta16-phi21*/	1, 21, 1, 
/* out0437_had-eta17-phi21*/	1, 21, 1, 
/* out0438_had-eta18-phi21*/	1, 21, 1, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 163, 5, 
/* out0442_had-eta2-phi22*/	3, 103, 1, 162, 1, 163, 3, 
/* out0443_had-eta3-phi22*/	4, 102, 3, 103, 10, 105, 2, 162, 5, 
/* out0444_had-eta4-phi22*/	4, 71, 1, 102, 10, 161, 2, 162, 2, 
/* out0445_had-eta5-phi22*/	4, 70, 1, 71, 4, 101, 4, 161, 4, 
/* out0446_had-eta6-phi22*/	3, 70, 7, 160, 2, 161, 2, 
/* out0447_had-eta7-phi22*/	4, 69, 3, 70, 3, 80, 1, 160, 3, 
/* out0448_had-eta8-phi22*/	3, 69, 5, 79, 1, 160, 2, 
/* out0449_had-eta9-phi22*/	4, 68, 1, 79, 4, 159, 3, 160, 1, 
/* out0450_had-eta10-phi22*/	4, 20, 1, 68, 1, 79, 2, 159, 5, 
/* out0451_had-eta11-phi22*/	1, 20, 3, 
/* out0452_had-eta12-phi22*/	1, 20, 3, 
/* out0453_had-eta13-phi22*/	3, 19, 1, 20, 1, 22, 1, 
/* out0454_had-eta14-phi22*/	2, 19, 1, 22, 1, 
/* out0455_had-eta15-phi22*/	2, 19, 1, 21, 1, 
/* out0456_had-eta16-phi22*/	1, 21, 1, 
/* out0457_had-eta17-phi22*/	1, 21, 1, 
/* out0458_had-eta18-phi22*/	1, 21, 1, 
/* out0459_had-eta19-phi22*/	1, 21, 1, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 168, 5, 
/* out0462_had-eta2-phi23*/	4, 73, 1, 103, 1, 167, 1, 168, 3, 
/* out0463_had-eta3-phi23*/	4, 72, 6, 73, 9, 103, 4, 167, 5, 
/* out0464_had-eta4-phi23*/	5, 71, 3, 72, 8, 82, 1, 166, 2, 167, 2, 
/* out0465_had-eta5-phi23*/	3, 71, 8, 81, 1, 166, 4, 
/* out0466_had-eta6-phi23*/	4, 70, 3, 81, 4, 165, 2, 166, 2, 
/* out0467_had-eta7-phi23*/	3, 70, 1, 80, 5, 165, 3, 
/* out0468_had-eta8-phi23*/	3, 79, 1, 80, 4, 165, 2, 
/* out0469_had-eta9-phi23*/	3, 79, 4, 164, 3, 165, 1, 
/* out0470_had-eta10-phi23*/	3, 23, 1, 79, 3, 164, 5, 
/* out0471_had-eta11-phi23*/	2, 20, 2, 23, 1, 
/* out0472_had-eta12-phi23*/	2, 20, 1, 22, 1, 
/* out0473_had-eta13-phi23*/	1, 22, 2, 
/* out0474_had-eta14-phi23*/	1, 22, 2, 
/* out0475_had-eta15-phi23*/	2, 21, 1, 22, 1, 
/* out0476_had-eta16-phi23*/	1, 21, 1, 
/* out0477_had-eta17-phi23*/	1, 21, 1, 
/* out0478_had-eta18-phi23*/	1, 21, 1, 
/* out0479_had-eta19-phi23*/	1, 21, 1, 
/* out0480_had-eta0-phi24*/	0, 
/* out0481_had-eta1-phi24*/	1, 168, 5, 
/* out0482_had-eta2-phi24*/	2, 167, 1, 168, 3, 
/* out0483_had-eta3-phi24*/	4, 72, 1, 73, 6, 83, 8, 167, 5, 
/* out0484_had-eta4-phi24*/	5, 72, 1, 82, 7, 83, 3, 166, 2, 167, 2, 
/* out0485_had-eta5-phi24*/	4, 81, 3, 82, 6, 91, 1, 166, 4, 
/* out0486_had-eta6-phi24*/	4, 81, 7, 90, 1, 165, 2, 166, 2, 
/* out0487_had-eta7-phi24*/	4, 80, 3, 81, 1, 90, 2, 165, 3, 
/* out0488_had-eta8-phi24*/	3, 80, 3, 89, 3, 165, 2, 
/* out0489_had-eta9-phi24*/	4, 79, 1, 89, 3, 164, 3, 165, 1, 
/* out0490_had-eta10-phi24*/	2, 23, 3, 164, 5, 
/* out0491_had-eta11-phi24*/	1, 23, 3, 
/* out0492_had-eta12-phi24*/	2, 22, 1, 23, 2, 
/* out0493_had-eta13-phi24*/	1, 22, 2, 
/* out0494_had-eta14-phi24*/	1, 22, 2, 
/* out0495_had-eta15-phi24*/	1, 22, 1, 
/* out0496_had-eta16-phi24*/	1, 21, 1, 
/* out0497_had-eta17-phi24*/	1, 21, 1, 
/* out0498_had-eta18-phi24*/	1, 21, 1, 
/* out0499_had-eta19-phi24*/	0, 
/* out0500_had-eta0-phi25*/	0, 
/* out0501_had-eta1-phi25*/	1, 173, 5, 
/* out0502_had-eta2-phi25*/	3, 93, 1, 172, 1, 173, 3, 
/* out0503_had-eta3-phi25*/	4, 83, 4, 92, 1, 93, 8, 172, 5, 
/* out0504_had-eta4-phi25*/	5, 82, 1, 83, 1, 92, 9, 171, 2, 172, 2, 
/* out0505_had-eta5-phi25*/	4, 82, 1, 91, 7, 92, 1, 171, 4, 
/* out0506_had-eta6-phi25*/	4, 90, 3, 91, 4, 170, 2, 171, 2, 
/* out0507_had-eta7-phi25*/	2, 90, 6, 170, 3, 
/* out0508_had-eta8-phi25*/	3, 89, 4, 90, 1, 170, 2, 
/* out0509_had-eta9-phi25*/	3, 89, 4, 169, 3, 170, 1, 
/* out0510_had-eta10-phi25*/	3, 23, 2, 89, 1, 169, 5, 
/* out0511_had-eta11-phi25*/	1, 23, 3, 
/* out0512_had-eta12-phi25*/	1, 23, 1, 
/* out0513_had-eta13-phi25*/	1, 22, 1, 
/* out0514_had-eta14-phi25*/	1, 22, 1, 
/* out0515_had-eta15-phi25*/	0, 
/* out0516_had-eta16-phi25*/	0, 
/* out0517_had-eta17-phi25*/	0, 
/* out0518_had-eta18-phi25*/	0, 
/* out0519_had-eta19-phi25*/	0, 
/* out0520_had-eta0-phi26*/	0, 
/* out0521_had-eta1-phi26*/	1, 173, 5, 
/* out0522_had-eta2-phi26*/	3, 93, 1, 172, 1, 173, 3, 
/* out0523_had-eta3-phi26*/	2, 93, 6, 172, 5, 
/* out0524_had-eta4-phi26*/	3, 92, 5, 171, 2, 172, 2, 
/* out0525_had-eta5-phi26*/	2, 91, 3, 171, 4, 
/* out0526_had-eta6-phi26*/	4, 90, 1, 91, 1, 170, 2, 171, 2, 
/* out0527_had-eta7-phi26*/	2, 90, 2, 170, 3, 
/* out0528_had-eta8-phi26*/	1, 170, 2, 
/* out0529_had-eta9-phi26*/	3, 89, 1, 169, 3, 170, 1, 
/* out0530_had-eta10-phi26*/	1, 169, 5, 
/* out0531_had-eta11-phi26*/	0, 
/* out0532_had-eta12-phi26*/	0, 
/* out0533_had-eta13-phi26*/	0, 
/* out0534_had-eta14-phi26*/	0, 
/* out0535_had-eta15-phi26*/	0, 
/* out0536_had-eta16-phi26*/	0, 
/* out0537_had-eta17-phi26*/	0, 
/* out0538_had-eta18-phi26*/	0, 
/* out0539_had-eta19-phi26*/	0, 
/* out0540_had-eta0-phi27*/	0, 
/* out0541_had-eta1-phi27*/	0, 
/* out0542_had-eta2-phi27*/	0, 
/* out0543_had-eta3-phi27*/	0, 
/* out0544_had-eta4-phi27*/	0, 
/* out0545_had-eta5-phi27*/	0, 
/* out0546_had-eta6-phi27*/	0, 
/* out0547_had-eta7-phi27*/	0, 
/* out0548_had-eta8-phi27*/	0, 
/* out0549_had-eta9-phi27*/	0, 
/* out0550_had-eta10-phi27*/	0, 
/* out0551_had-eta11-phi27*/	0, 
/* out0552_had-eta12-phi27*/	0, 
/* out0553_had-eta13-phi27*/	0, 
/* out0554_had-eta14-phi27*/	0, 
/* out0555_had-eta15-phi27*/	0, 
/* out0556_had-eta16-phi27*/	0, 
/* out0557_had-eta17-phi27*/	0, 
/* out0558_had-eta18-phi27*/	0, 
/* out0559_had-eta19-phi27*/	0, 
};