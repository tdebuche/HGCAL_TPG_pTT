parameter integer matrixE [0:1904] = {
/* num inputs = 108(in0-in107) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 3 */
//* total number of input in adders 672 */

/* out0000_em-eta0-phi0*/	0, 
/* out0001_em-eta1-phi0*/	0, 
/* out0002_em-eta2-phi0*/	0, 
/* out0003_em-eta3-phi0*/	0, 
/* out0004_em-eta4-phi0*/	0, 
/* out0005_em-eta5-phi0*/	0, 
/* out0006_em-eta6-phi0*/	0, 
/* out0007_em-eta7-phi0*/	0, 
/* out0008_em-eta8-phi0*/	0, 
/* out0009_em-eta9-phi0*/	0, 
/* out0010_em-eta10-phi0*/	0, 
/* out0011_em-eta11-phi0*/	0, 
/* out0012_em-eta12-phi0*/	0, 
/* out0013_em-eta13-phi0*/	0, 
/* out0014_em-eta14-phi0*/	0, 
/* out0015_em-eta15-phi0*/	0, 
/* out0016_em-eta16-phi0*/	0, 
/* out0017_em-eta17-phi0*/	0, 
/* out0018_em-eta18-phi0*/	0, 
/* out0019_em-eta19-phi0*/	1, 0, 1, 
/* out0020_em-eta0-phi1*/	0, 
/* out0021_em-eta1-phi1*/	0, 
/* out0022_em-eta2-phi1*/	0, 
/* out0023_em-eta3-phi1*/	0, 
/* out0024_em-eta4-phi1*/	0, 
/* out0025_em-eta5-phi1*/	0, 
/* out0026_em-eta6-phi1*/	0, 
/* out0027_em-eta7-phi1*/	0, 
/* out0028_em-eta8-phi1*/	0, 
/* out0029_em-eta9-phi1*/	0, 
/* out0030_em-eta10-phi1*/	0, 
/* out0031_em-eta11-phi1*/	0, 
/* out0032_em-eta12-phi1*/	1, 2, 1, 
/* out0033_em-eta13-phi1*/	0, 
/* out0034_em-eta14-phi1*/	1, 1, 1, 
/* out0035_em-eta15-phi1*/	1, 1, 1, 
/* out0036_em-eta16-phi1*/	1, 1, 1, 
/* out0037_em-eta17-phi1*/	1, 0, 1, 
/* out0038_em-eta18-phi1*/	1, 0, 1, 
/* out0039_em-eta19-phi1*/	1, 0, 1, 
/* out0040_em-eta0-phi2*/	0, 
/* out0041_em-eta1-phi2*/	0, 
/* out0042_em-eta2-phi2*/	0, 
/* out0043_em-eta3-phi2*/	1, 41, 8, 
/* out0044_em-eta4-phi2*/	1, 40, 6, 
/* out0045_em-eta5-phi2*/	2, 39, 3, 40, 1, 
/* out0046_em-eta6-phi2*/	1, 39, 4, 
/* out0047_em-eta7-phi2*/	1, 38, 5, 
/* out0048_em-eta8-phi2*/	2, 37, 1, 38, 3, 
/* out0049_em-eta9-phi2*/	1, 37, 4, 
/* out0050_em-eta10-phi2*/	1, 37, 3, 
/* out0051_em-eta11-phi2*/	1, 2, 3, 
/* out0052_em-eta12-phi2*/	1, 2, 2, 
/* out0053_em-eta13-phi2*/	1, 2, 1, 
/* out0054_em-eta14-phi2*/	1, 1, 2, 
/* out0055_em-eta15-phi2*/	1, 1, 1, 
/* out0056_em-eta16-phi2*/	1, 1, 1, 
/* out0057_em-eta17-phi2*/	2, 0, 1, 1, 1, 
/* out0058_em-eta18-phi2*/	1, 0, 1, 
/* out0059_em-eta19-phi2*/	1, 0, 1, 
/* out0060_em-eta0-phi3*/	0, 
/* out0061_em-eta1-phi3*/	0, 
/* out0062_em-eta2-phi3*/	1, 36, 3, 
/* out0063_em-eta3-phi3*/	3, 35, 3, 36, 4, 41, 8, 
/* out0064_em-eta4-phi3*/	3, 34, 1, 35, 2, 40, 7, 
/* out0065_em-eta5-phi3*/	3, 34, 3, 39, 4, 40, 2, 
/* out0066_em-eta6-phi3*/	2, 33, 2, 39, 5, 
/* out0067_em-eta7-phi3*/	1, 38, 5, 
/* out0068_em-eta8-phi3*/	3, 32, 1, 37, 1, 38, 3, 
/* out0069_em-eta9-phi3*/	1, 37, 4, 
/* out0070_em-eta10-phi3*/	1, 37, 3, 
/* out0071_em-eta11-phi3*/	1, 2, 3, 
/* out0072_em-eta12-phi3*/	1, 2, 2, 
/* out0073_em-eta13-phi3*/	1, 2, 2, 
/* out0074_em-eta14-phi3*/	1, 1, 2, 
/* out0075_em-eta15-phi3*/	1, 1, 1, 
/* out0076_em-eta16-phi3*/	1, 1, 1, 
/* out0077_em-eta17-phi3*/	2, 0, 1, 1, 1, 
/* out0078_em-eta18-phi3*/	1, 0, 2, 
/* out0079_em-eta19-phi3*/	1, 0, 1, 
/* out0080_em-eta0-phi4*/	0, 
/* out0081_em-eta1-phi4*/	0, 
/* out0082_em-eta2-phi4*/	2, 31, 1, 36, 4, 
/* out0083_em-eta3-phi4*/	3, 31, 4, 35, 6, 36, 5, 
/* out0084_em-eta4-phi4*/	3, 30, 2, 34, 3, 35, 5, 
/* out0085_em-eta5-phi4*/	1, 34, 8, 
/* out0086_em-eta6-phi4*/	1, 33, 7, 
/* out0087_em-eta7-phi4*/	2, 32, 2, 33, 4, 
/* out0088_em-eta8-phi4*/	1, 32, 5, 
/* out0089_em-eta9-phi4*/	2, 6, 1, 32, 2, 
/* out0090_em-eta10-phi4*/	1, 6, 3, 
/* out0091_em-eta11-phi4*/	2, 2, 1, 6, 2, 
/* out0092_em-eta12-phi4*/	2, 2, 1, 5, 1, 
/* out0093_em-eta13-phi4*/	1, 5, 2, 
/* out0094_em-eta14-phi4*/	2, 1, 1, 5, 1, 
/* out0095_em-eta15-phi4*/	1, 1, 1, 
/* out0096_em-eta16-phi4*/	1, 1, 1, 
/* out0097_em-eta17-phi4*/	1, 0, 1, 
/* out0098_em-eta18-phi4*/	1, 0, 1, 
/* out0099_em-eta19-phi4*/	1, 0, 1, 
/* out0100_em-eta0-phi5*/	0, 
/* out0101_em-eta1-phi5*/	0, 
/* out0102_em-eta2-phi5*/	1, 31, 3, 
/* out0103_em-eta3-phi5*/	3, 30, 2, 31, 8, 45, 2, 
/* out0104_em-eta4-phi5*/	1, 30, 10, 
/* out0105_em-eta5-phi5*/	3, 29, 7, 30, 1, 34, 1, 
/* out0106_em-eta6-phi5*/	3, 28, 1, 29, 3, 33, 2, 
/* out0107_em-eta7-phi5*/	3, 28, 4, 32, 1, 33, 1, 
/* out0108_em-eta8-phi5*/	1, 32, 4, 
/* out0109_em-eta9-phi5*/	3, 6, 2, 27, 1, 32, 1, 
/* out0110_em-eta10-phi5*/	1, 6, 3, 
/* out0111_em-eta11-phi5*/	1, 6, 3, 
/* out0112_em-eta12-phi5*/	1, 5, 2, 
/* out0113_em-eta13-phi5*/	1, 5, 2, 
/* out0114_em-eta14-phi5*/	1, 5, 2, 
/* out0115_em-eta15-phi5*/	1, 4, 1, 
/* out0116_em-eta16-phi5*/	1, 4, 1, 
/* out0117_em-eta17-phi5*/	1, 4, 1, 
/* out0118_em-eta18-phi5*/	2, 0, 1, 4, 1, 
/* out0119_em-eta19-phi5*/	1, 0, 1, 
/* out0120_em-eta0-phi6*/	0, 
/* out0121_em-eta1-phi6*/	0, 
/* out0122_em-eta2-phi6*/	2, 45, 1, 53, 4, 
/* out0123_em-eta3-phi6*/	2, 45, 12, 53, 1, 
/* out0124_em-eta4-phi6*/	3, 30, 1, 44, 8, 45, 1, 
/* out0125_em-eta5-phi6*/	3, 29, 4, 43, 2, 44, 3, 
/* out0126_em-eta6-phi6*/	3, 28, 3, 29, 2, 43, 2, 
/* out0127_em-eta7-phi6*/	1, 28, 6, 
/* out0128_em-eta8-phi6*/	2, 27, 4, 28, 1, 
/* out0129_em-eta9-phi6*/	1, 27, 4, 
/* out0130_em-eta10-phi6*/	3, 6, 1, 11, 1, 27, 1, 
/* out0131_em-eta11-phi6*/	2, 6, 1, 11, 2, 
/* out0132_em-eta12-phi6*/	1, 5, 2, 
/* out0133_em-eta13-phi6*/	1, 5, 2, 
/* out0134_em-eta14-phi6*/	1, 5, 1, 
/* out0135_em-eta15-phi6*/	1, 4, 1, 
/* out0136_em-eta16-phi6*/	1, 4, 1, 
/* out0137_em-eta17-phi6*/	1, 4, 1, 
/* out0138_em-eta18-phi6*/	1, 4, 1, 
/* out0139_em-eta19-phi6*/	1, 3, 1, 
/* out0140_em-eta0-phi7*/	0, 
/* out0141_em-eta1-phi7*/	0, 
/* out0142_em-eta2-phi7*/	1, 53, 7, 
/* out0143_em-eta3-phi7*/	2, 51, 9, 53, 4, 
/* out0144_em-eta4-phi7*/	3, 44, 4, 50, 2, 51, 3, 
/* out0145_em-eta5-phi7*/	3, 43, 5, 44, 1, 50, 2, 
/* out0146_em-eta6-phi7*/	2, 42, 1, 43, 6, 
/* out0147_em-eta7-phi7*/	2, 28, 1, 42, 5, 
/* out0148_em-eta8-phi7*/	2, 27, 3, 42, 2, 
/* out0149_em-eta9-phi7*/	1, 27, 3, 
/* out0150_em-eta10-phi7*/	1, 11, 3, 
/* out0151_em-eta11-phi7*/	1, 11, 3, 
/* out0152_em-eta12-phi7*/	1, 11, 1, 
/* out0153_em-eta13-phi7*/	2, 5, 1, 10, 1, 
/* out0154_em-eta14-phi7*/	1, 10, 1, 
/* out0155_em-eta15-phi7*/	1, 4, 1, 
/* out0156_em-eta16-phi7*/	1, 4, 1, 
/* out0157_em-eta17-phi7*/	1, 4, 1, 
/* out0158_em-eta18-phi7*/	2, 3, 1, 4, 1, 
/* out0159_em-eta19-phi7*/	1, 3, 2, 
/* out0160_em-eta0-phi8*/	0, 
/* out0161_em-eta1-phi8*/	0, 
/* out0162_em-eta2-phi8*/	0, 
/* out0163_em-eta3-phi8*/	2, 51, 3, 52, 6, 
/* out0164_em-eta4-phi8*/	3, 50, 7, 51, 1, 52, 2, 
/* out0165_em-eta5-phi8*/	2, 46, 3, 50, 5, 
/* out0166_em-eta6-phi8*/	3, 42, 1, 43, 1, 46, 5, 
/* out0167_em-eta7-phi8*/	1, 42, 5, 
/* out0168_em-eta8-phi8*/	2, 22, 3, 42, 2, 
/* out0169_em-eta9-phi8*/	1, 22, 4, 
/* out0170_em-eta10-phi8*/	2, 11, 2, 22, 1, 
/* out0171_em-eta11-phi8*/	1, 11, 3, 
/* out0172_em-eta12-phi8*/	2, 10, 1, 11, 1, 
/* out0173_em-eta13-phi8*/	1, 10, 2, 
/* out0174_em-eta14-phi8*/	1, 10, 2, 
/* out0175_em-eta15-phi8*/	2, 4, 1, 10, 1, 
/* out0176_em-eta16-phi8*/	1, 4, 1, 
/* out0177_em-eta17-phi8*/	1, 4, 1, 
/* out0178_em-eta18-phi8*/	2, 3, 1, 4, 1, 
/* out0179_em-eta19-phi8*/	1, 3, 3, 
/* out0180_em-eta0-phi9*/	0, 
/* out0181_em-eta1-phi9*/	0, 
/* out0182_em-eta2-phi9*/	0, 
/* out0183_em-eta3-phi9*/	2, 48, 3, 52, 6, 
/* out0184_em-eta4-phi9*/	3, 47, 7, 48, 1, 52, 2, 
/* out0185_em-eta5-phi9*/	2, 46, 3, 47, 5, 
/* out0186_em-eta6-phi9*/	3, 23, 1, 24, 1, 46, 5, 
/* out0187_em-eta7-phi9*/	1, 23, 5, 
/* out0188_em-eta8-phi9*/	2, 22, 3, 23, 2, 
/* out0189_em-eta9-phi9*/	1, 22, 4, 
/* out0190_em-eta10-phi9*/	2, 12, 2, 22, 1, 
/* out0191_em-eta11-phi9*/	1, 12, 2, 
/* out0192_em-eta12-phi9*/	2, 10, 1, 12, 1, 
/* out0193_em-eta13-phi9*/	1, 10, 2, 
/* out0194_em-eta14-phi9*/	1, 10, 2, 
/* out0195_em-eta15-phi9*/	2, 7, 1, 10, 1, 
/* out0196_em-eta16-phi9*/	1, 7, 1, 
/* out0197_em-eta17-phi9*/	1, 7, 1, 
/* out0198_em-eta18-phi9*/	2, 3, 1, 7, 1, 
/* out0199_em-eta19-phi9*/	1, 3, 3, 
/* out0200_em-eta0-phi10*/	0, 
/* out0201_em-eta1-phi10*/	0, 
/* out0202_em-eta2-phi10*/	1, 49, 7, 
/* out0203_em-eta3-phi10*/	2, 48, 9, 49, 4, 
/* out0204_em-eta4-phi10*/	3, 25, 4, 47, 2, 48, 3, 
/* out0205_em-eta5-phi10*/	3, 24, 5, 25, 1, 47, 2, 
/* out0206_em-eta6-phi10*/	2, 23, 1, 24, 6, 
/* out0207_em-eta7-phi10*/	2, 18, 1, 23, 5, 
/* out0208_em-eta8-phi10*/	2, 17, 3, 23, 2, 
/* out0209_em-eta9-phi10*/	1, 17, 3, 
/* out0210_em-eta10-phi10*/	1, 12, 3, 
/* out0211_em-eta11-phi10*/	1, 12, 3, 
/* out0212_em-eta12-phi10*/	1, 12, 2, 
/* out0213_em-eta13-phi10*/	2, 8, 1, 10, 1, 
/* out0214_em-eta14-phi10*/	1, 10, 1, 
/* out0215_em-eta15-phi10*/	1, 7, 1, 
/* out0216_em-eta16-phi10*/	1, 7, 1, 
/* out0217_em-eta17-phi10*/	1, 7, 1, 
/* out0218_em-eta18-phi10*/	2, 3, 1, 7, 1, 
/* out0219_em-eta19-phi10*/	1, 3, 2, 
/* out0220_em-eta0-phi11*/	0, 
/* out0221_em-eta1-phi11*/	0, 
/* out0222_em-eta2-phi11*/	2, 26, 1, 49, 4, 
/* out0223_em-eta3-phi11*/	2, 26, 12, 49, 1, 
/* out0224_em-eta4-phi11*/	3, 20, 1, 25, 8, 26, 1, 
/* out0225_em-eta5-phi11*/	3, 19, 4, 24, 2, 25, 3, 
/* out0226_em-eta6-phi11*/	3, 18, 3, 19, 2, 24, 2, 
/* out0227_em-eta7-phi11*/	1, 18, 6, 
/* out0228_em-eta8-phi11*/	2, 17, 4, 18, 1, 
/* out0229_em-eta9-phi11*/	1, 17, 4, 
/* out0230_em-eta10-phi11*/	3, 9, 1, 12, 1, 17, 1, 
/* out0231_em-eta11-phi11*/	2, 9, 1, 12, 2, 
/* out0232_em-eta12-phi11*/	1, 8, 2, 
/* out0233_em-eta13-phi11*/	1, 8, 2, 
/* out0234_em-eta14-phi11*/	1, 8, 1, 
/* out0235_em-eta15-phi11*/	1, 7, 1, 
/* out0236_em-eta16-phi11*/	1, 7, 1, 
/* out0237_em-eta17-phi11*/	1, 7, 1, 
/* out0238_em-eta18-phi11*/	1, 7, 1, 
/* out0239_em-eta19-phi11*/	1, 3, 1, 
/* out0240_em-eta0-phi12*/	0, 
/* out0241_em-eta1-phi12*/	0, 
/* out0242_em-eta2-phi12*/	1, 21, 3, 
/* out0243_em-eta3-phi12*/	3, 20, 2, 21, 8, 26, 2, 
/* out0244_em-eta4-phi12*/	1, 20, 10, 
/* out0245_em-eta5-phi12*/	3, 15, 1, 19, 7, 20, 1, 
/* out0246_em-eta6-phi12*/	3, 14, 2, 18, 1, 19, 3, 
/* out0247_em-eta7-phi12*/	3, 13, 1, 14, 1, 18, 4, 
/* out0248_em-eta8-phi12*/	1, 13, 4, 
/* out0249_em-eta9-phi12*/	3, 9, 2, 13, 1, 17, 1, 
/* out0250_em-eta10-phi12*/	1, 9, 3, 
/* out0251_em-eta11-phi12*/	1, 9, 3, 
/* out0252_em-eta12-phi12*/	1, 8, 2, 
/* out0253_em-eta13-phi12*/	1, 8, 2, 
/* out0254_em-eta14-phi12*/	1, 8, 2, 
/* out0255_em-eta15-phi12*/	1, 7, 1, 
/* out0256_em-eta16-phi12*/	1, 7, 1, 
/* out0257_em-eta17-phi12*/	1, 7, 1, 
/* out0258_em-eta18-phi12*/	1, 7, 1, 
/* out0259_em-eta19-phi12*/	1, 54, 1, 
/* out0260_em-eta0-phi13*/	0, 
/* out0261_em-eta1-phi13*/	0, 
/* out0262_em-eta2-phi13*/	1, 21, 1, 
/* out0263_em-eta3-phi13*/	2, 16, 6, 21, 4, 
/* out0264_em-eta4-phi13*/	3, 15, 3, 16, 5, 20, 2, 
/* out0265_em-eta5-phi13*/	1, 15, 8, 
/* out0266_em-eta6-phi13*/	1, 14, 7, 
/* out0267_em-eta7-phi13*/	2, 13, 2, 14, 4, 
/* out0268_em-eta8-phi13*/	1, 13, 5, 
/* out0269_em-eta9-phi13*/	2, 9, 1, 13, 2, 
/* out0270_em-eta10-phi13*/	1, 9, 3, 
/* out0271_em-eta11-phi13*/	1, 9, 2, 
/* out0272_em-eta12-phi13*/	2, 8, 1, 56, 1, 
/* out0273_em-eta13-phi13*/	1, 8, 2, 
/* out0274_em-eta14-phi13*/	2, 8, 1, 55, 1, 
/* out0275_em-eta15-phi13*/	1, 55, 1, 
/* out0276_em-eta16-phi13*/	1, 55, 1, 
/* out0277_em-eta17-phi13*/	1, 54, 1, 
/* out0278_em-eta18-phi13*/	1, 54, 1, 
/* out0279_em-eta19-phi13*/	1, 54, 1, 
/* out0280_em-eta0-phi14*/	0, 
/* out0281_em-eta1-phi14*/	0, 
/* out0282_em-eta2-phi14*/	0, 
/* out0283_em-eta3-phi14*/	2, 16, 3, 95, 8, 
/* out0284_em-eta4-phi14*/	3, 15, 1, 16, 2, 94, 6, 
/* out0285_em-eta5-phi14*/	3, 15, 3, 93, 3, 94, 1, 
/* out0286_em-eta6-phi14*/	2, 14, 2, 93, 4, 
/* out0287_em-eta7-phi14*/	1, 92, 5, 
/* out0288_em-eta8-phi14*/	3, 13, 1, 91, 1, 92, 3, 
/* out0289_em-eta9-phi14*/	1, 91, 4, 
/* out0290_em-eta10-phi14*/	1, 91, 3, 
/* out0291_em-eta11-phi14*/	1, 56, 3, 
/* out0292_em-eta12-phi14*/	1, 56, 2, 
/* out0293_em-eta13-phi14*/	1, 56, 1, 
/* out0294_em-eta14-phi14*/	1, 55, 2, 
/* out0295_em-eta15-phi14*/	1, 55, 1, 
/* out0296_em-eta16-phi14*/	1, 55, 1, 
/* out0297_em-eta17-phi14*/	2, 54, 1, 55, 1, 
/* out0298_em-eta18-phi14*/	1, 54, 1, 
/* out0299_em-eta19-phi14*/	1, 54, 1, 
/* out0300_em-eta0-phi15*/	0, 
/* out0301_em-eta1-phi15*/	0, 
/* out0302_em-eta2-phi15*/	1, 90, 3, 
/* out0303_em-eta3-phi15*/	3, 89, 3, 90, 4, 95, 8, 
/* out0304_em-eta4-phi15*/	3, 88, 1, 89, 2, 94, 7, 
/* out0305_em-eta5-phi15*/	3, 88, 3, 93, 4, 94, 2, 
/* out0306_em-eta6-phi15*/	2, 87, 2, 93, 5, 
/* out0307_em-eta7-phi15*/	1, 92, 5, 
/* out0308_em-eta8-phi15*/	3, 86, 1, 91, 1, 92, 3, 
/* out0309_em-eta9-phi15*/	1, 91, 4, 
/* out0310_em-eta10-phi15*/	1, 91, 3, 
/* out0311_em-eta11-phi15*/	1, 56, 3, 
/* out0312_em-eta12-phi15*/	1, 56, 2, 
/* out0313_em-eta13-phi15*/	1, 56, 2, 
/* out0314_em-eta14-phi15*/	1, 55, 2, 
/* out0315_em-eta15-phi15*/	1, 55, 1, 
/* out0316_em-eta16-phi15*/	1, 55, 1, 
/* out0317_em-eta17-phi15*/	2, 54, 1, 55, 1, 
/* out0318_em-eta18-phi15*/	1, 54, 2, 
/* out0319_em-eta19-phi15*/	1, 54, 1, 
/* out0320_em-eta0-phi16*/	0, 
/* out0321_em-eta1-phi16*/	0, 
/* out0322_em-eta2-phi16*/	2, 85, 1, 90, 4, 
/* out0323_em-eta3-phi16*/	3, 85, 4, 89, 6, 90, 5, 
/* out0324_em-eta4-phi16*/	3, 84, 2, 88, 3, 89, 5, 
/* out0325_em-eta5-phi16*/	1, 88, 8, 
/* out0326_em-eta6-phi16*/	1, 87, 7, 
/* out0327_em-eta7-phi16*/	2, 86, 2, 87, 4, 
/* out0328_em-eta8-phi16*/	1, 86, 5, 
/* out0329_em-eta9-phi16*/	2, 60, 1, 86, 2, 
/* out0330_em-eta10-phi16*/	1, 60, 3, 
/* out0331_em-eta11-phi16*/	2, 56, 1, 60, 2, 
/* out0332_em-eta12-phi16*/	2, 56, 1, 59, 1, 
/* out0333_em-eta13-phi16*/	1, 59, 2, 
/* out0334_em-eta14-phi16*/	2, 55, 1, 59, 1, 
/* out0335_em-eta15-phi16*/	1, 55, 1, 
/* out0336_em-eta16-phi16*/	1, 55, 1, 
/* out0337_em-eta17-phi16*/	1, 54, 1, 
/* out0338_em-eta18-phi16*/	1, 54, 1, 
/* out0339_em-eta19-phi16*/	1, 54, 1, 
/* out0340_em-eta0-phi17*/	0, 
/* out0341_em-eta1-phi17*/	0, 
/* out0342_em-eta2-phi17*/	1, 85, 3, 
/* out0343_em-eta3-phi17*/	3, 84, 2, 85, 8, 99, 2, 
/* out0344_em-eta4-phi17*/	1, 84, 10, 
/* out0345_em-eta5-phi17*/	3, 83, 7, 84, 1, 88, 1, 
/* out0346_em-eta6-phi17*/	3, 82, 1, 83, 3, 87, 2, 
/* out0347_em-eta7-phi17*/	3, 82, 4, 86, 1, 87, 1, 
/* out0348_em-eta8-phi17*/	1, 86, 4, 
/* out0349_em-eta9-phi17*/	3, 60, 2, 81, 1, 86, 1, 
/* out0350_em-eta10-phi17*/	1, 60, 3, 
/* out0351_em-eta11-phi17*/	1, 60, 3, 
/* out0352_em-eta12-phi17*/	1, 59, 2, 
/* out0353_em-eta13-phi17*/	1, 59, 2, 
/* out0354_em-eta14-phi17*/	1, 59, 2, 
/* out0355_em-eta15-phi17*/	1, 58, 1, 
/* out0356_em-eta16-phi17*/	1, 58, 1, 
/* out0357_em-eta17-phi17*/	1, 58, 1, 
/* out0358_em-eta18-phi17*/	2, 54, 1, 58, 1, 
/* out0359_em-eta19-phi17*/	1, 54, 1, 
/* out0360_em-eta0-phi18*/	0, 
/* out0361_em-eta1-phi18*/	0, 
/* out0362_em-eta2-phi18*/	2, 99, 1, 107, 4, 
/* out0363_em-eta3-phi18*/	2, 99, 12, 107, 1, 
/* out0364_em-eta4-phi18*/	3, 84, 1, 98, 8, 99, 1, 
/* out0365_em-eta5-phi18*/	3, 83, 4, 97, 2, 98, 3, 
/* out0366_em-eta6-phi18*/	3, 82, 3, 83, 2, 97, 2, 
/* out0367_em-eta7-phi18*/	1, 82, 6, 
/* out0368_em-eta8-phi18*/	2, 81, 4, 82, 1, 
/* out0369_em-eta9-phi18*/	1, 81, 4, 
/* out0370_em-eta10-phi18*/	3, 60, 1, 66, 1, 81, 1, 
/* out0371_em-eta11-phi18*/	2, 60, 1, 66, 2, 
/* out0372_em-eta12-phi18*/	1, 59, 2, 
/* out0373_em-eta13-phi18*/	1, 59, 2, 
/* out0374_em-eta14-phi18*/	1, 59, 1, 
/* out0375_em-eta15-phi18*/	1, 58, 1, 
/* out0376_em-eta16-phi18*/	1, 58, 1, 
/* out0377_em-eta17-phi18*/	1, 58, 1, 
/* out0378_em-eta18-phi18*/	1, 58, 1, 
/* out0379_em-eta19-phi18*/	1, 57, 1, 
/* out0380_em-eta0-phi19*/	0, 
/* out0381_em-eta1-phi19*/	0, 
/* out0382_em-eta2-phi19*/	1, 107, 7, 
/* out0383_em-eta3-phi19*/	2, 106, 9, 107, 4, 
/* out0384_em-eta4-phi19*/	3, 98, 4, 104, 2, 106, 3, 
/* out0385_em-eta5-phi19*/	3, 97, 5, 98, 1, 104, 2, 
/* out0386_em-eta6-phi19*/	2, 96, 1, 97, 6, 
/* out0387_em-eta7-phi19*/	2, 82, 1, 96, 5, 
/* out0388_em-eta8-phi19*/	2, 81, 3, 96, 2, 
/* out0389_em-eta9-phi19*/	1, 81, 3, 
/* out0390_em-eta10-phi19*/	1, 66, 3, 
/* out0391_em-eta11-phi19*/	1, 66, 3, 
/* out0392_em-eta12-phi19*/	1, 66, 1, 
/* out0393_em-eta13-phi19*/	2, 59, 1, 64, 1, 
/* out0394_em-eta14-phi19*/	1, 64, 1, 
/* out0395_em-eta15-phi19*/	1, 58, 1, 
/* out0396_em-eta16-phi19*/	1, 58, 1, 
/* out0397_em-eta17-phi19*/	1, 58, 1, 
/* out0398_em-eta18-phi19*/	2, 57, 1, 58, 1, 
/* out0399_em-eta19-phi19*/	1, 57, 2, 
/* out0400_em-eta0-phi20*/	0, 
/* out0401_em-eta1-phi20*/	0, 
/* out0402_em-eta2-phi20*/	0, 
/* out0403_em-eta3-phi20*/	2, 105, 6, 106, 3, 
/* out0404_em-eta4-phi20*/	3, 104, 7, 105, 2, 106, 1, 
/* out0405_em-eta5-phi20*/	2, 100, 3, 104, 5, 
/* out0406_em-eta6-phi20*/	3, 96, 1, 97, 1, 100, 5, 
/* out0407_em-eta7-phi20*/	1, 96, 5, 
/* out0408_em-eta8-phi20*/	2, 76, 3, 96, 2, 
/* out0409_em-eta9-phi20*/	1, 76, 4, 
/* out0410_em-eta10-phi20*/	2, 66, 2, 76, 1, 
/* out0411_em-eta11-phi20*/	1, 66, 3, 
/* out0412_em-eta12-phi20*/	2, 64, 1, 66, 1, 
/* out0413_em-eta13-phi20*/	1, 64, 2, 
/* out0414_em-eta14-phi20*/	1, 64, 2, 
/* out0415_em-eta15-phi20*/	2, 58, 1, 64, 1, 
/* out0416_em-eta16-phi20*/	1, 58, 1, 
/* out0417_em-eta17-phi20*/	1, 58, 1, 
/* out0418_em-eta18-phi20*/	2, 57, 1, 58, 1, 
/* out0419_em-eta19-phi20*/	1, 57, 3, 
/* out0420_em-eta0-phi21*/	0, 
/* out0421_em-eta1-phi21*/	0, 
/* out0422_em-eta2-phi21*/	0, 
/* out0423_em-eta3-phi21*/	2, 102, 3, 105, 6, 
/* out0424_em-eta4-phi21*/	3, 101, 7, 102, 1, 105, 2, 
/* out0425_em-eta5-phi21*/	2, 100, 3, 101, 5, 
/* out0426_em-eta6-phi21*/	3, 77, 1, 78, 1, 100, 5, 
/* out0427_em-eta7-phi21*/	1, 77, 5, 
/* out0428_em-eta8-phi21*/	2, 76, 3, 77, 2, 
/* out0429_em-eta9-phi21*/	1, 76, 4, 
/* out0430_em-eta10-phi21*/	2, 65, 2, 76, 1, 
/* out0431_em-eta11-phi21*/	1, 65, 2, 
/* out0432_em-eta12-phi21*/	2, 64, 1, 65, 1, 
/* out0433_em-eta13-phi21*/	1, 64, 2, 
/* out0434_em-eta14-phi21*/	1, 64, 2, 
/* out0435_em-eta15-phi21*/	2, 61, 1, 64, 1, 
/* out0436_em-eta16-phi21*/	1, 61, 1, 
/* out0437_em-eta17-phi21*/	1, 61, 1, 
/* out0438_em-eta18-phi21*/	2, 57, 1, 61, 1, 
/* out0439_em-eta19-phi21*/	1, 57, 3, 
/* out0440_em-eta0-phi22*/	0, 
/* out0441_em-eta1-phi22*/	0, 
/* out0442_em-eta2-phi22*/	1, 103, 7, 
/* out0443_em-eta3-phi22*/	2, 102, 9, 103, 4, 
/* out0444_em-eta4-phi22*/	3, 79, 4, 101, 2, 102, 3, 
/* out0445_em-eta5-phi22*/	3, 78, 5, 79, 1, 101, 2, 
/* out0446_em-eta6-phi22*/	2, 77, 1, 78, 6, 
/* out0447_em-eta7-phi22*/	2, 72, 1, 77, 5, 
/* out0448_em-eta8-phi22*/	2, 71, 3, 77, 2, 
/* out0449_em-eta9-phi22*/	1, 71, 3, 
/* out0450_em-eta10-phi22*/	1, 65, 3, 
/* out0451_em-eta11-phi22*/	1, 65, 3, 
/* out0452_em-eta12-phi22*/	1, 65, 2, 
/* out0453_em-eta13-phi22*/	2, 62, 1, 64, 1, 
/* out0454_em-eta14-phi22*/	1, 64, 1, 
/* out0455_em-eta15-phi22*/	1, 61, 1, 
/* out0456_em-eta16-phi22*/	1, 61, 1, 
/* out0457_em-eta17-phi22*/	1, 61, 1, 
/* out0458_em-eta18-phi22*/	2, 57, 1, 61, 1, 
/* out0459_em-eta19-phi22*/	1, 57, 2, 
/* out0460_em-eta0-phi23*/	0, 
/* out0461_em-eta1-phi23*/	0, 
/* out0462_em-eta2-phi23*/	2, 80, 1, 103, 4, 
/* out0463_em-eta3-phi23*/	2, 80, 12, 103, 1, 
/* out0464_em-eta4-phi23*/	3, 74, 1, 79, 8, 80, 1, 
/* out0465_em-eta5-phi23*/	3, 73, 4, 78, 2, 79, 3, 
/* out0466_em-eta6-phi23*/	3, 72, 3, 73, 2, 78, 2, 
/* out0467_em-eta7-phi23*/	1, 72, 6, 
/* out0468_em-eta8-phi23*/	2, 71, 4, 72, 1, 
/* out0469_em-eta9-phi23*/	1, 71, 4, 
/* out0470_em-eta10-phi23*/	3, 63, 1, 65, 1, 71, 1, 
/* out0471_em-eta11-phi23*/	2, 63, 1, 65, 2, 
/* out0472_em-eta12-phi23*/	1, 62, 2, 
/* out0473_em-eta13-phi23*/	1, 62, 2, 
/* out0474_em-eta14-phi23*/	1, 62, 1, 
/* out0475_em-eta15-phi23*/	1, 61, 1, 
/* out0476_em-eta16-phi23*/	1, 61, 1, 
/* out0477_em-eta17-phi23*/	1, 61, 1, 
/* out0478_em-eta18-phi23*/	1, 61, 1, 
/* out0479_em-eta19-phi23*/	1, 57, 1, 
/* out0480_em-eta0-phi24*/	0, 
/* out0481_em-eta1-phi24*/	0, 
/* out0482_em-eta2-phi24*/	1, 75, 3, 
/* out0483_em-eta3-phi24*/	3, 74, 2, 75, 8, 80, 2, 
/* out0484_em-eta4-phi24*/	1, 74, 10, 
/* out0485_em-eta5-phi24*/	3, 69, 1, 73, 7, 74, 1, 
/* out0486_em-eta6-phi24*/	3, 68, 2, 72, 1, 73, 3, 
/* out0487_em-eta7-phi24*/	3, 67, 1, 68, 1, 72, 4, 
/* out0488_em-eta8-phi24*/	1, 67, 4, 
/* out0489_em-eta9-phi24*/	3, 63, 2, 67, 1, 71, 1, 
/* out0490_em-eta10-phi24*/	1, 63, 3, 
/* out0491_em-eta11-phi24*/	1, 63, 3, 
/* out0492_em-eta12-phi24*/	1, 62, 2, 
/* out0493_em-eta13-phi24*/	1, 62, 2, 
/* out0494_em-eta14-phi24*/	1, 62, 2, 
/* out0495_em-eta15-phi24*/	1, 61, 1, 
/* out0496_em-eta16-phi24*/	1, 61, 1, 
/* out0497_em-eta17-phi24*/	1, 61, 1, 
/* out0498_em-eta18-phi24*/	1, 61, 1, 
/* out0499_em-eta19-phi24*/	0, 
/* out0500_em-eta0-phi25*/	0, 
/* out0501_em-eta1-phi25*/	0, 
/* out0502_em-eta2-phi25*/	1, 75, 1, 
/* out0503_em-eta3-phi25*/	2, 70, 6, 75, 4, 
/* out0504_em-eta4-phi25*/	3, 69, 3, 70, 5, 74, 2, 
/* out0505_em-eta5-phi25*/	1, 69, 8, 
/* out0506_em-eta6-phi25*/	1, 68, 7, 
/* out0507_em-eta7-phi25*/	2, 67, 2, 68, 4, 
/* out0508_em-eta8-phi25*/	1, 67, 5, 
/* out0509_em-eta9-phi25*/	2, 63, 1, 67, 2, 
/* out0510_em-eta10-phi25*/	1, 63, 3, 
/* out0511_em-eta11-phi25*/	1, 63, 2, 
/* out0512_em-eta12-phi25*/	1, 62, 1, 
/* out0513_em-eta13-phi25*/	1, 62, 2, 
/* out0514_em-eta14-phi25*/	1, 62, 1, 
/* out0515_em-eta15-phi25*/	0, 
/* out0516_em-eta16-phi25*/	0, 
/* out0517_em-eta17-phi25*/	0, 
/* out0518_em-eta18-phi25*/	0, 
/* out0519_em-eta19-phi25*/	0, 
/* out0520_em-eta0-phi26*/	0, 
/* out0521_em-eta1-phi26*/	0, 
/* out0522_em-eta2-phi26*/	0, 
/* out0523_em-eta3-phi26*/	1, 70, 3, 
/* out0524_em-eta4-phi26*/	2, 69, 1, 70, 2, 
/* out0525_em-eta5-phi26*/	1, 69, 3, 
/* out0526_em-eta6-phi26*/	1, 68, 2, 
/* out0527_em-eta7-phi26*/	0, 
/* out0528_em-eta8-phi26*/	1, 67, 1, 
/* out0529_em-eta9-phi26*/	0, 
/* out0530_em-eta10-phi26*/	0, 
/* out0531_em-eta11-phi26*/	0, 
/* out0532_em-eta12-phi26*/	0, 
/* out0533_em-eta13-phi26*/	0, 
/* out0534_em-eta14-phi26*/	0, 
/* out0535_em-eta15-phi26*/	0, 
/* out0536_em-eta16-phi26*/	0, 
/* out0537_em-eta17-phi26*/	0, 
/* out0538_em-eta18-phi26*/	0, 
/* out0539_em-eta19-phi26*/	0, 
/* out0540_em-eta0-phi27*/	0, 
/* out0541_em-eta1-phi27*/	0, 
/* out0542_em-eta2-phi27*/	0, 
/* out0543_em-eta3-phi27*/	0, 
/* out0544_em-eta4-phi27*/	0, 
/* out0545_em-eta5-phi27*/	0, 
/* out0546_em-eta6-phi27*/	0, 
/* out0547_em-eta7-phi27*/	0, 
/* out0548_em-eta8-phi27*/	0, 
/* out0549_em-eta9-phi27*/	0, 
/* out0550_em-eta10-phi27*/	0, 
/* out0551_em-eta11-phi27*/	0, 
/* out0552_em-eta12-phi27*/	0, 
/* out0553_em-eta13-phi27*/	0, 
/* out0554_em-eta14-phi27*/	0, 
/* out0555_em-eta15-phi27*/	0, 
/* out0556_em-eta16-phi27*/	0, 
/* out0557_em-eta17-phi27*/	0, 
/* out0558_em-eta18-phi27*/	0, 
/* out0559_em-eta19-phi27*/	0, 
};