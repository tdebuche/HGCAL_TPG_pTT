parameter integer matrixH [0:4409] = {
/* num inputs = 112(in0-in111) */
/* num outputs = 600(out0-out599) */
//* max inputs per outputs = 11 */
//* total number of input in adders 1269 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	0,
/* out0006_em-eta6-phi0*/	0,
/* out0007_em-eta7-phi0*/	0,
/* out0008_em-eta8-phi0*/	0,
/* out0009_em-eta9-phi0*/	0,
/* out0010_em-eta10-phi0*/	0,
/* out0011_em-eta11-phi0*/	0,
/* out0012_em-eta12-phi0*/	0,
/* out0013_em-eta13-phi0*/	0,
/* out0014_em-eta14-phi0*/	0,
/* out0015_em-eta15-phi0*/	0,
/* out0016_em-eta16-phi0*/	0,
/* out0017_em-eta17-phi0*/	0,
/* out0018_em-eta18-phi0*/	0,
/* out0019_em-eta19-phi0*/	0,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	0,
/* out0026_em-eta6-phi1*/	0,
/* out0027_em-eta7-phi1*/	0,
/* out0028_em-eta8-phi1*/	0,
/* out0029_em-eta9-phi1*/	0,
/* out0030_em-eta10-phi1*/	0,
/* out0031_em-eta11-phi1*/	0,
/* out0032_em-eta12-phi1*/	0,
/* out0033_em-eta13-phi1*/	0,
/* out0034_em-eta14-phi1*/	0,
/* out0035_em-eta15-phi1*/	0,
/* out0036_em-eta16-phi1*/	0,
/* out0037_em-eta17-phi1*/	0,
/* out0038_em-eta18-phi1*/	0,
/* out0039_em-eta19-phi1*/	0,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	0,
/* out0046_em-eta6-phi2*/	0,
/* out0047_em-eta7-phi2*/	0,
/* out0048_em-eta8-phi2*/	0,
/* out0049_em-eta9-phi2*/	0,
/* out0050_em-eta10-phi2*/	0,
/* out0051_em-eta11-phi2*/	0,
/* out0052_em-eta12-phi2*/	0,
/* out0053_em-eta13-phi2*/	0,
/* out0054_em-eta14-phi2*/	0,
/* out0055_em-eta15-phi2*/	0,
/* out0056_em-eta16-phi2*/	0,
/* out0057_em-eta17-phi2*/	0,
/* out0058_em-eta18-phi2*/	0,
/* out0059_em-eta19-phi2*/	0,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	0,
/* out0065_em-eta5-phi3*/	0,
/* out0066_em-eta6-phi3*/	0,
/* out0067_em-eta7-phi3*/	0,
/* out0068_em-eta8-phi3*/	0,
/* out0069_em-eta9-phi3*/	2,42,0,4,42,2,1,
/* out0070_em-eta10-phi3*/	1,42,2,3,
/* out0071_em-eta11-phi3*/	2,33,0,4,33,2,1,
/* out0072_em-eta12-phi3*/	1,33,2,3,
/* out0073_em-eta13-phi3*/	1,24,0,4,
/* out0074_em-eta14-phi3*/	1,24,2,4,
/* out0075_em-eta15-phi3*/	1,15,0,1,
/* out0076_em-eta16-phi3*/	1,15,0,3,
/* out0077_em-eta17-phi3*/	1,15,2,3,
/* out0078_em-eta18-phi3*/	1,15,2,1,
/* out0079_em-eta19-phi3*/	0,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	0,
/* out0085_em-eta5-phi4*/	0,
/* out0086_em-eta6-phi4*/	0,
/* out0087_em-eta7-phi4*/	0,
/* out0088_em-eta8-phi4*/	0,
/* out0089_em-eta9-phi4*/	5,42,0,12,42,1,5,42,2,1,101,1,3,101,2,13,
/* out0090_em-eta10-phi4*/	6,33,0,3,42,1,2,42,2,11,93,0,8,93,1,3,101,1,1,
/* out0091_em-eta11-phi4*/	5,33,0,9,33,1,3,33,2,2,93,0,8,93,2,2,
/* out0092_em-eta12-phi4*/	5,24,0,1,33,1,1,33,2,9,85,0,7,85,1,1,
/* out0093_em-eta13-phi4*/	3,24,0,9,24,1,1,85,0,7,
/* out0094_em-eta14-phi4*/	4,24,1,1,24,2,7,77,0,2,77,1,1,
/* out0095_em-eta15-phi4*/	3,15,0,4,24,2,3,77,0,6,
/* out0096_em-eta16-phi4*/	2,15,0,5,77,0,3,
/* out0097_em-eta17-phi4*/	2,15,2,5,70,2,2,
/* out0098_em-eta18-phi4*/	3,15,2,3,70,0,1,70,2,3,
/* out0099_em-eta19-phi4*/	0,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	0,
/* out0105_em-eta5-phi5*/	0,
/* out0106_em-eta6-phi5*/	0,
/* out0107_em-eta7-phi5*/	0,
/* out0108_em-eta8-phi5*/	0,
/* out0109_em-eta9-phi5*/	7,42,1,5,43,0,2,50,1,4,50,2,13,101,1,11,101,2,3,102,0,5,
/* out0110_em-eta10-phi5*/	7,42,1,4,43,0,9,43,2,3,93,1,13,93,2,1,101,1,1,102,0,3,
/* out0111_em-eta11-phi5*/	6,33,1,8,34,0,1,43,2,5,85,1,1,93,2,12,94,0,1,
/* out0112_em-eta12-phi5*/	7,24,0,1,33,1,4,33,2,1,34,0,5,34,2,1,85,0,1,85,1,11,
/* out0113_em-eta13-phi5*/	5,24,0,1,24,1,7,34,2,2,85,0,1,85,2,9,
/* out0114_em-eta14-phi5*/	4,24,1,7,24,2,1,77,1,6,85,2,2,
/* out0115_em-eta15-phi5*/	7,15,0,2,15,1,2,24,2,1,25,2,1,77,0,4,77,1,2,77,2,2,
/* out0116_em-eta16-phi5*/	4,15,0,1,15,1,5,77,0,1,77,2,4,
/* out0117_em-eta17-phi5*/	3,15,1,3,15,2,2,70,2,6,
/* out0118_em-eta18-phi5*/	3,15,2,2,70,0,3,70,2,2,
/* out0119_em-eta19-phi5*/	0,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	0,
/* out0125_em-eta5-phi6*/	0,
/* out0126_em-eta6-phi6*/	0,
/* out0127_em-eta7-phi6*/	0,
/* out0128_em-eta8-phi6*/	3,50,1,1,50,2,2,51,0,1,
/* out0129_em-eta9-phi6*/	11,43,0,2,43,1,1,50,1,11,50,2,1,51,0,11,51,2,3,102,0,4,102,1,13,102,2,2,108,0,1,108,1,1,
/* out0130_em-eta10-phi6*/	7,43,0,3,43,1,11,43,2,2,93,2,1,94,1,3,102,0,4,102,2,9,
/* out0131_em-eta11-phi6*/	7,34,0,5,34,1,1,43,1,2,43,2,6,94,0,10,94,1,4,94,2,1,
/* out0132_em-eta12-phi6*/	8,34,0,5,34,1,3,34,2,3,85,1,3,85,2,1,86,1,1,94,0,5,94,2,2,
/* out0133_em-eta13-phi6*/	4,25,0,2,34,2,8,85,2,4,86,0,6,
/* out0134_em-eta14-phi6*/	3,25,0,8,77,1,5,86,0,4,
/* out0135_em-eta15-phi6*/	4,25,0,1,25,2,6,77,1,2,77,2,4,
/* out0136_em-eta16-phi6*/	6,15,1,3,16,1,1,25,2,2,70,2,1,77,2,5,78,0,1,
/* out0137_em-eta17-phi6*/	4,15,1,2,16,1,2,70,0,4,70,2,2,
/* out0138_em-eta18-phi6*/	3,15,1,1,16,1,2,70,0,3,
/* out0139_em-eta19-phi6*/	0,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	0,
/* out0145_em-eta5-phi7*/	0,
/* out0146_em-eta6-phi7*/	0,
/* out0147_em-eta7-phi7*/	0,
/* out0148_em-eta8-phi7*/	1,51,1,1,
/* out0149_em-eta9-phi7*/	10,51,0,4,51,1,10,51,2,7,102,1,3,102,2,2,103,0,2,103,1,4,108,0,14,108,1,14,108,2,14,
/* out0150_em-eta10-phi7*/	6,43,1,2,44,0,10,51,2,5,94,1,3,102,2,3,103,0,11,
/* out0151_em-eta11-phi7*/	6,34,1,2,44,0,4,44,2,8,94,1,6,94,2,7,103,0,1,
/* out0152_em-eta12-phi7*/	6,34,1,8,35,0,2,44,2,1,86,1,5,94,2,6,95,0,1,
/* out0153_em-eta13-phi7*/	9,25,0,2,25,1,2,34,1,2,34,2,2,35,0,2,35,2,1,86,0,3,86,1,6,86,2,2,
/* out0154_em-eta14-phi7*/	4,25,0,3,25,1,5,86,0,3,86,2,5,
/* out0155_em-eta15-phi7*/	5,25,1,2,25,2,5,77,2,1,78,0,3,78,1,2,
/* out0156_em-eta16-phi7*/	3,16,2,3,25,2,2,78,0,6,
/* out0157_em-eta17-phi7*/	4,16,1,3,16,2,1,70,0,3,78,0,2,
/* out0158_em-eta18-phi7*/	2,16,1,3,70,0,2,
/* out0159_em-eta19-phi7*/	0,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	0,
/* out0165_em-eta5-phi8*/	0,
/* out0166_em-eta6-phi8*/	0,
/* out0167_em-eta7-phi8*/	0,
/* out0168_em-eta8-phi8*/	0,
/* out0169_em-eta9-phi8*/	11,51,1,5,52,0,16,52,1,3,52,2,2,103,1,10,108,0,1,108,1,1,108,2,2,109,0,8,109,1,5,109,2,3,
/* out0170_em-eta10-phi8*/	7,44,0,2,44,1,9,51,2,1,52,2,5,103,0,2,103,1,2,103,2,13,
/* out0171_em-eta11-phi8*/	5,44,1,7,44,2,6,95,0,5,95,1,8,103,2,2,
/* out0172_em-eta12-phi8*/	6,35,0,10,35,1,1,44,2,1,86,1,1,95,0,10,95,2,1,
/* out0173_em-eta13-phi8*/	5,35,0,2,35,2,8,86,1,3,86,2,4,87,0,1,
/* out0174_em-eta14-phi8*/	6,25,1,4,26,0,2,35,2,2,78,1,2,86,2,5,87,0,2,
/* out0175_em-eta15-phi8*/	3,25,1,3,26,0,3,78,1,7,
/* out0176_em-eta16-phi8*/	5,16,2,5,26,2,1,78,0,2,78,1,1,78,2,3,
/* out0177_em-eta17-phi8*/	5,16,0,1,16,1,1,16,2,3,78,0,2,78,2,3,
/* out0178_em-eta18-phi8*/	1,16,1,3,
/* out0179_em-eta19-phi8*/	0,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	0,
/* out0185_em-eta5-phi9*/	0,
/* out0186_em-eta6-phi9*/	0,
/* out0187_em-eta7-phi9*/	0,
/* out0188_em-eta8-phi9*/	0,
/* out0189_em-eta9-phi9*/	6,52,1,12,52,2,1,104,1,6,109,0,8,109,1,11,109,2,13,
/* out0190_em-eta10-phi9*/	6,45,0,8,52,1,1,52,2,8,103,2,1,104,0,13,104,1,2,
/* out0191_em-eta11-phi9*/	5,45,0,8,45,2,6,95,1,8,95,2,4,104,0,3,
/* out0192_em-eta12-phi9*/	4,35,1,10,45,2,2,87,1,1,95,2,11,
/* out0193_em-eta13-phi9*/	4,35,1,5,35,2,4,87,0,3,87,1,7,
/* out0194_em-eta14-phi9*/	3,26,0,7,35,2,1,87,0,8,
/* out0195_em-eta15-phi9*/	5,26,0,4,26,2,3,78,1,4,78,2,2,87,0,2,
/* out0196_em-eta16-phi9*/	3,16,2,2,26,2,4,78,2,6,
/* out0197_em-eta17-phi9*/	3,16,0,8,16,2,2,78,2,2,
/* out0198_em-eta18-phi9*/	2,16,0,7,16,1,1,
/* out0199_em-eta19-phi9*/	0,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	0,
/* out0205_em-eta5-phi10*/	0,
/* out0206_em-eta6-phi10*/	0,
/* out0207_em-eta7-phi10*/	0,
/* out0208_em-eta8-phi10*/	0,
/* out0209_em-eta9-phi10*/	7,53,0,15,53,1,6,53,2,2,104,1,6,110,0,13,110,1,11,110,2,8,
/* out0210_em-eta10-phi10*/	6,45,1,8,53,0,1,53,2,8,104,1,2,104,2,13,105,0,1,
/* out0211_em-eta11-phi10*/	5,45,1,8,45,2,6,96,0,4,96,1,8,104,2,3,
/* out0212_em-eta12-phi10*/	4,36,0,10,45,2,2,87,1,1,96,0,11,
/* out0213_em-eta13-phi10*/	4,36,0,5,36,2,4,87,1,7,87,2,3,
/* out0214_em-eta14-phi10*/	3,26,1,7,36,2,1,87,2,8,
/* out0215_em-eta15-phi10*/	5,26,1,4,26,2,3,79,0,2,79,1,4,87,2,2,
/* out0216_em-eta16-phi10*/	3,17,2,1,26,2,4,79,0,6,
/* out0217_em-eta17-phi10*/	3,17,1,3,17,2,1,79,0,2,
/* out0218_em-eta18-phi10*/	1,17,1,3,
/* out0219_em-eta19-phi10*/	0,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	0,
/* out0225_em-eta5-phi11*/	0,
/* out0226_em-eta6-phi11*/	0,
/* out0227_em-eta7-phi11*/	0,
/* out0228_em-eta8-phi11*/	0,
/* out0229_em-eta9-phi11*/	11,53,1,10,53,2,1,54,0,10,54,1,1,105,1,10,110,0,3,110,1,5,110,2,8,111,0,2,111,1,1,111,2,1,
/* out0230_em-eta10-phi11*/	6,46,0,9,46,1,2,53,2,5,105,0,13,105,1,2,105,2,2,
/* out0231_em-eta11-phi11*/	5,46,0,7,46,2,6,96,1,8,96,2,5,105,0,2,
/* out0232_em-eta12-phi11*/	6,36,0,1,36,1,10,46,2,1,88,1,1,96,0,1,96,2,10,
/* out0233_em-eta13-phi11*/	5,36,1,2,36,2,8,87,2,1,88,0,4,88,1,3,
/* out0234_em-eta14-phi11*/	6,26,1,2,27,0,4,36,2,2,79,1,2,87,2,2,88,0,5,
/* out0235_em-eta15-phi11*/	3,26,1,3,27,0,3,79,1,7,
/* out0236_em-eta16-phi11*/	5,17,2,5,26,2,1,79,0,3,79,1,1,79,2,2,
/* out0237_em-eta17-phi11*/	4,17,1,2,17,2,3,79,0,3,79,2,2,
/* out0238_em-eta18-phi11*/	1,17,1,3,
/* out0239_em-eta19-phi11*/	0,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	0,
/* out0245_em-eta5-phi12*/	0,
/* out0246_em-eta6-phi12*/	0,
/* out0247_em-eta7-phi12*/	0,
/* out0248_em-eta8-phi12*/	1,54,1,1,
/* out0249_em-eta9-phi12*/	10,54,0,6,54,1,9,54,2,8,105,1,4,105,2,2,106,0,2,106,1,3,111,0,14,111,1,14,111,2,14,
/* out0250_em-eta10-phi12*/	6,46,1,10,47,0,2,54,2,5,97,1,3,105,2,11,106,0,3,
/* out0251_em-eta11-phi12*/	6,37,0,2,46,1,4,46,2,8,97,0,7,97,1,6,105,2,1,
/* out0252_em-eta12-phi12*/	6,36,1,2,37,0,8,46,2,1,88,1,5,96,2,1,97,0,6,
/* out0253_em-eta13-phi12*/	9,27,0,2,27,1,2,36,1,2,36,2,1,37,0,2,37,2,2,88,0,2,88,1,6,88,2,3,
/* out0254_em-eta14-phi12*/	4,27,0,5,27,1,3,88,0,5,88,2,3,
/* out0255_em-eta15-phi12*/	5,27,0,2,27,2,5,79,1,2,79,2,3,80,0,1,
/* out0256_em-eta16-phi12*/	3,17,2,4,27,2,2,79,2,6,
/* out0257_em-eta17-phi12*/	5,17,0,7,17,1,1,17,2,2,71,1,3,79,2,2,
/* out0258_em-eta18-phi12*/	2,17,1,3,71,1,2,
/* out0259_em-eta19-phi12*/	0,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	0,
/* out0265_em-eta5-phi13*/	0,
/* out0266_em-eta6-phi13*/	0,
/* out0267_em-eta7-phi13*/	0,
/* out0268_em-eta8-phi13*/	2,54,1,1,55,0,3,
/* out0269_em-eta9-phi13*/	11,47,0,1,47,1,2,54,1,4,54,2,3,55,0,9,55,2,3,106,0,2,106,1,13,106,2,4,111,1,1,111,2,1,
/* out0270_em-eta10-phi13*/	7,47,0,11,47,1,3,47,2,2,97,1,3,98,0,1,106,0,9,106,2,4,
/* out0271_em-eta11-phi13*/	7,37,0,1,37,1,5,47,0,2,47,2,6,97,0,1,97,1,4,97,2,10,
/* out0272_em-eta12-phi13*/	8,37,0,3,37,1,5,37,2,3,88,1,1,89,0,1,89,1,3,97,0,2,97,2,5,
/* out0273_em-eta13-phi13*/	4,27,1,2,37,2,8,88,2,6,89,0,4,
/* out0274_em-eta14-phi13*/	3,27,1,8,80,1,5,88,2,4,
/* out0275_em-eta15-phi13*/	4,27,1,1,27,2,6,80,0,4,80,1,2,
/* out0276_em-eta16-phi13*/	6,17,0,1,18,0,3,27,2,2,71,2,1,79,2,1,80,0,5,
/* out0277_em-eta17-phi13*/	4,17,0,6,18,0,2,71,1,4,71,2,2,
/* out0278_em-eta18-phi13*/	4,17,0,2,17,1,1,18,0,1,71,1,3,
/* out0279_em-eta19-phi13*/	0,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	0,
/* out0285_em-eta5-phi14*/	0,
/* out0286_em-eta6-phi14*/	0,
/* out0287_em-eta7-phi14*/	0,
/* out0288_em-eta8-phi14*/	0,
/* out0289_em-eta9-phi14*/	7,47,1,2,48,0,5,55,0,4,55,2,13,106,2,5,107,0,12,107,2,3,
/* out0290_em-eta10-phi14*/	7,47,1,9,47,2,3,48,0,4,98,0,1,98,1,13,106,2,3,107,2,1,
/* out0291_em-eta11-phi14*/	6,37,1,1,38,0,8,47,2,5,89,1,1,97,2,1,98,0,12,
/* out0292_em-eta12-phi14*/	7,28,1,1,37,1,5,37,2,1,38,0,4,38,2,1,89,1,11,89,2,1,
/* out0293_em-eta13-phi14*/	5,28,0,7,28,1,1,37,2,2,89,0,9,89,2,1,
/* out0294_em-eta14-phi14*/	4,28,0,7,28,2,1,80,1,6,89,0,2,
/* out0295_em-eta15-phi14*/	7,18,0,2,18,1,2,27,2,1,28,2,1,80,0,2,80,1,2,80,2,4,
/* out0296_em-eta16-phi14*/	4,18,0,5,18,1,1,80,0,4,80,2,1,
/* out0297_em-eta17-phi14*/	3,18,0,3,18,2,2,71,2,6,
/* out0298_em-eta18-phi14*/	3,18,2,2,71,1,3,71,2,2,
/* out0299_em-eta19-phi14*/	0,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	0,
/* out0305_em-eta5-phi15*/	0,
/* out0306_em-eta6-phi15*/	0,
/* out0307_em-eta7-phi15*/	0,
/* out0308_em-eta8-phi15*/	0,
/* out0309_em-eta9-phi15*/	6,48,0,5,48,1,12,48,2,1,99,1,3,107,0,4,107,2,11,
/* out0310_em-eta10-phi15*/	8,38,1,3,48,0,2,48,2,11,98,1,3,98,2,8,99,0,4,99,1,1,107,2,1,
/* out0311_em-eta11-phi15*/	6,38,0,3,38,1,9,38,2,2,90,1,4,98,0,2,98,2,8,
/* out0312_em-eta12-phi15*/	6,28,1,1,38,0,1,38,2,9,89,1,1,89,2,7,90,0,4,
/* out0313_em-eta13-phi15*/	4,28,0,1,28,1,9,81,1,2,89,2,7,
/* out0314_em-eta14-phi15*/	6,28,0,1,28,2,7,80,1,1,80,2,2,81,0,3,81,1,2,
/* out0315_em-eta15-phi15*/	4,18,1,4,28,2,3,80,2,6,81,0,1,
/* out0316_em-eta16-phi15*/	3,18,1,5,72,1,3,80,2,3,
/* out0317_em-eta17-phi15*/	3,18,2,5,71,2,2,72,0,3,
/* out0318_em-eta18-phi15*/	4,18,2,3,71,1,1,71,2,3,72,0,1,
/* out0319_em-eta19-phi15*/	0,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	0,
/* out0325_em-eta5-phi16*/	0,
/* out0326_em-eta6-phi16*/	0,
/* out0327_em-eta7-phi16*/	0,
/* out0328_em-eta8-phi16*/	0,
/* out0329_em-eta9-phi16*/	7,39,1,1,48,1,4,48,2,1,49,0,13,49,2,4,99,1,11,99,2,4,
/* out0330_em-eta10-phi16*/	6,39,0,11,39,1,3,48,2,3,99,0,12,99,1,1,99,2,4,
/* out0331_em-eta11-phi16*/	7,29,1,1,38,1,4,38,2,1,39,0,5,39,2,2,90,1,12,90,2,2,
/* out0332_em-eta12-phi16*/	5,29,0,8,29,1,1,38,2,3,90,0,10,90,2,1,
/* out0333_em-eta13-phi16*/	4,28,1,4,29,0,6,81,1,9,90,0,1,
/* out0334_em-eta14-phi16*/	6,19,0,3,19,1,1,28,2,4,81,0,6,81,1,2,81,2,1,
/* out0335_em-eta15-phi16*/	4,18,1,1,19,0,6,72,1,3,81,0,4,
/* out0336_em-eta16-phi16*/	3,18,1,3,19,0,2,72,1,6,
/* out0337_em-eta17-phi16*/	4,9,1,2,18,2,3,72,0,4,72,1,1,
/* out0338_em-eta18-phi16*/	3,9,1,3,18,2,1,72,0,4,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	0,
/* out0345_em-eta5-phi17*/	0,
/* out0346_em-eta6-phi17*/	0,
/* out0347_em-eta7-phi17*/	0,
/* out0348_em-eta8-phi17*/	0,
/* out0349_em-eta9-phi17*/	7,39,1,1,40,0,6,49,0,3,49,2,12,99,2,3,100,0,13,100,2,4,
/* out0350_em-eta10-phi17*/	6,39,1,11,39,2,4,40,0,1,91,0,1,91,1,10,99,2,5,
/* out0351_em-eta11-phi17*/	6,29,1,3,30,0,1,39,2,9,82,1,1,90,2,7,91,0,7,
/* out0352_em-eta12-phi17*/	6,29,0,1,29,1,8,29,2,2,82,1,5,90,0,1,90,2,6,
/* out0353_em-eta13-phi17*/	5,29,0,1,29,2,9,81,1,1,81,2,6,82,0,3,
/* out0354_em-eta14-phi17*/	3,19,0,1,19,1,7,81,2,8,
/* out0355_em-eta15-phi17*/	9,19,0,3,19,1,1,19,2,2,72,1,2,72,2,1,73,0,1,73,1,1,81,0,2,81,2,1,
/* out0356_em-eta16-phi17*/	5,9,2,1,19,0,1,19,2,4,72,1,1,72,2,4,
/* out0357_em-eta17-phi17*/	4,9,1,4,9,2,3,72,0,1,72,2,4,
/* out0358_em-eta18-phi17*/	2,9,1,3,72,0,3,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	0,
/* out0365_em-eta5-phi18*/	0,
/* out0366_em-eta6-phi18*/	0,
/* out0367_em-eta7-phi18*/	0,
/* out0368_em-eta8-phi18*/	3,40,1,3,41,0,1,41,1,1,
/* out0369_em-eta9-phi18*/	8,40,0,6,40,1,10,40,2,4,91,1,1,92,0,13,92,2,2,100,0,3,100,2,12,
/* out0370_em-eta10-phi18*/	9,30,0,1,30,1,5,39,2,1,40,0,3,40,2,6,91,0,1,91,1,5,91,2,11,92,2,1,
/* out0371_em-eta11-phi18*/	7,30,0,11,30,1,2,30,2,1,82,1,3,82,2,1,91,0,7,91,2,3,
/* out0372_em-eta12-phi18*/	9,20,0,1,20,1,1,29,1,3,29,2,2,30,0,3,30,2,2,82,0,1,82,1,7,82,2,3,
/* out0373_em-eta13-phi18*/	3,20,0,7,29,2,3,82,0,10,
/* out0374_em-eta14-phi18*/	3,19,1,6,20,0,2,73,1,8,
/* out0375_em-eta15-phi18*/	4,19,1,1,19,2,6,73,0,4,73,1,3,
/* out0376_em-eta16-phi18*/	5,9,2,2,10,0,1,19,2,3,72,2,3,73,0,3,
/* out0377_em-eta17-phi18*/	4,9,1,1,9,2,6,65,1,2,72,2,3,
/* out0378_em-eta18-phi18*/	3,9,1,2,65,1,2,72,2,1,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	0,
/* out0385_em-eta5-phi19*/	0,
/* out0386_em-eta6-phi19*/	0,
/* out0387_em-eta7-phi19*/	0,
/* out0388_em-eta8-phi19*/	3,41,0,3,41,1,1,41,2,3,
/* out0389_em-eta9-phi19*/	10,31,0,4,31,1,4,40,1,3,40,2,4,41,0,11,41,1,13,41,2,11,92,0,3,92,1,11,92,2,4,
/* out0390_em-eta10-phi19*/	6,30,1,5,31,0,10,40,2,2,83,1,7,91,2,2,92,2,9,
/* out0391_em-eta11-phi19*/	5,30,1,4,30,2,9,82,2,1,83,0,7,83,1,7,
/* out0392_em-eta12-phi19*/	6,20,1,7,21,0,1,30,2,4,74,1,2,82,2,8,83,0,2,
/* out0393_em-eta13-phi19*/	9,20,0,4,20,1,3,20,2,3,73,1,1,73,2,1,74,0,1,74,1,2,82,0,2,82,2,3,
/* out0394_em-eta14-phi19*/	5,10,1,1,20,0,2,20,2,4,73,1,3,73,2,5,
/* out0395_em-eta15-phi19*/	5,10,0,4,10,1,2,19,2,1,73,0,4,73,2,3,
/* out0396_em-eta16-phi19*/	3,10,0,6,65,2,2,73,0,3,
/* out0397_em-eta17-phi19*/	4,9,2,4,10,0,2,65,1,3,65,2,2,
/* out0398_em-eta18-phi19*/	2,9,1,1,65,1,3,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	0,
/* out0405_em-eta5-phi20*/	0,
/* out0406_em-eta6-phi20*/	0,
/* out0407_em-eta7-phi20*/	0,
/* out0408_em-eta8-phi20*/	0,
/* out0409_em-eta9-phi20*/	11,31,1,12,31,2,1,32,0,8,32,1,5,32,2,3,41,0,1,41,1,1,41,2,2,84,0,13,84,1,3,92,1,4,
/* out0410_em-eta10-phi20*/	8,21,1,2,31,0,2,31,2,13,83,1,2,83,2,7,84,0,3,84,2,7,92,1,1,
/* out0411_em-eta11-phi20*/	4,21,0,7,21,1,6,83,0,5,83,2,9,
/* out0412_em-eta12-phi20*/	6,20,1,3,21,0,8,21,2,1,74,1,8,74,2,1,83,0,2,
/* out0413_em-eta13-phi20*/	5,11,0,2,20,1,2,20,2,6,74,0,6,74,1,4,
/* out0414_em-eta14-phi20*/	6,10,1,3,11,0,1,20,2,3,66,1,1,73,2,3,74,0,4,
/* out0415_em-eta15-phi20*/	3,10,1,6,66,1,3,73,2,4,
/* out0416_em-eta16-phi20*/	6,10,0,2,10,2,3,65,2,4,66,0,1,66,1,1,73,0,1,
/* out0417_em-eta17-phi20*/	4,10,0,1,10,2,2,65,0,1,65,2,4,
/* out0418_em-eta18-phi20*/	2,65,0,1,65,1,3,
/* out0419_em-eta19-phi20*/	1,65,1,1,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	0,
/* out0425_em-eta5-phi21*/	0,
/* out0426_em-eta6-phi21*/	0,
/* out0427_em-eta7-phi21*/	0,
/* out0428_em-eta8-phi21*/	0,
/* out0429_em-eta9-phi21*/	7,22,0,2,22,1,7,31,2,1,32,0,8,32,1,11,32,2,13,84,1,10,
/* out0430_em-eta10-phi21*/	7,21,1,1,22,0,13,22,1,1,31,2,1,75,1,6,84,1,3,84,2,9,
/* out0431_em-eta11-phi21*/	5,21,1,7,21,2,6,22,0,1,75,0,4,75,1,10,
/* out0432_em-eta12-phi21*/	4,11,1,3,21,2,9,74,2,8,75,0,4,
/* out0433_em-eta13-phi21*/	4,11,0,5,11,1,5,74,0,3,74,2,7,
/* out0434_em-eta14-phi21*/	4,10,1,1,11,0,7,66,1,6,74,0,2,
/* out0435_em-eta15-phi21*/	5,10,1,3,10,2,3,11,0,1,66,0,2,66,1,5,
/* out0436_em-eta16-phi21*/	3,10,2,6,65,2,1,66,0,5,
/* out0437_em-eta17-phi21*/	3,10,2,2,65,0,5,65,2,3,
/* out0438_em-eta18-phi21*/	2,65,0,8,65,1,1,
/* out0439_em-eta19-phi21*/	2,65,0,1,65,1,1,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	0,
/* out0445_em-eta5-phi22*/	0,
/* out0446_em-eta6-phi22*/	0,
/* out0447_em-eta7-phi22*/	0,
/* out0448_em-eta8-phi22*/	0,
/* out0449_em-eta9-phi22*/	8,13,0,1,22,1,7,22,2,2,23,0,13,23,1,11,23,2,8,76,0,10,76,1,6,
/* out0450_em-eta10-phi22*/	7,12,1,1,13,0,1,22,1,1,22,2,13,75,2,6,76,0,6,76,2,10,
/* out0451_em-eta11-phi22*/	5,12,0,6,12,1,7,22,2,1,75,0,4,75,2,10,
/* out0452_em-eta12-phi22*/	4,11,1,3,12,0,9,67,1,8,75,0,4,
/* out0453_em-eta13-phi22*/	4,11,1,5,11,2,5,67,0,3,67,1,7,
/* out0454_em-eta14-phi22*/	4,5,1,1,11,2,7,66,2,6,67,0,2,
/* out0455_em-eta15-phi22*/	5,5,0,3,5,1,3,11,2,1,66,0,2,66,2,5,
/* out0456_em-eta16-phi22*/	3,5,0,6,60,2,1,66,0,5,
/* out0457_em-eta17-phi22*/	3,5,0,2,60,1,2,60,2,2,
/* out0458_em-eta18-phi22*/	1,60,1,3,
/* out0459_em-eta19-phi22*/	1,60,1,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	0,
/* out0465_em-eta5-phi23*/	0,
/* out0466_em-eta6-phi23*/	0,
/* out0467_em-eta7-phi23*/	0,
/* out0468_em-eta8-phi23*/	0,
/* out0469_em-eta9-phi23*/	11,13,0,1,13,1,12,14,0,2,14,1,1,14,2,1,23,0,3,23,1,5,23,2,8,69,0,8,69,1,1,76,1,8,
/* out0470_em-eta10-phi23*/	9,12,1,2,13,0,13,13,2,2,68,1,7,68,2,2,69,0,2,69,2,1,76,1,2,76,2,6,
/* out0471_em-eta11-phi23*/	4,12,1,6,12,2,7,68,0,5,68,1,9,
/* out0472_em-eta12-phi23*/	6,6,1,3,12,0,1,12,2,8,67,1,1,67,2,8,68,0,2,
/* out0473_em-eta13-phi23*/	5,6,0,6,6,1,2,11,2,2,67,0,6,67,2,4,
/* out0474_em-eta14-phi23*/	6,5,1,3,6,0,3,11,2,1,61,1,3,66,2,1,67,0,4,
/* out0475_em-eta15-phi23*/	3,5,1,6,61,1,4,66,2,3,
/* out0476_em-eta16-phi23*/	6,5,0,3,5,2,2,60,2,4,61,0,1,66,0,1,66,2,1,
/* out0477_em-eta17-phi23*/	4,5,0,2,5,2,1,60,1,1,60,2,4,
/* out0478_em-eta18-phi23*/	1,60,1,4,
/* out0479_em-eta19-phi23*/	1,60,1,1,
/* out0480_em-eta0-phi24*/	0,
/* out0481_em-eta1-phi24*/	0,
/* out0482_em-eta2-phi24*/	0,
/* out0483_em-eta3-phi24*/	0,
/* out0484_em-eta4-phi24*/	0,
/* out0485_em-eta5-phi24*/	0,
/* out0486_em-eta6-phi24*/	0,
/* out0487_em-eta7-phi24*/	0,
/* out0488_em-eta8-phi24*/	3,14,0,3,14,1,1,14,2,3,
/* out0489_em-eta9-phi24*/	10,8,0,4,8,1,3,13,1,4,13,2,4,14,0,11,14,1,13,14,2,11,69,0,6,69,1,10,69,2,4,
/* out0490_em-eta10-phi24*/	6,7,1,5,8,0,2,13,2,10,63,1,2,68,2,7,69,2,9,
/* out0491_em-eta11-phi24*/	5,7,0,9,7,1,4,62,1,1,68,0,7,68,2,7,
/* out0492_em-eta12-phi24*/	6,6,1,7,7,0,4,12,2,1,62,1,8,67,2,2,68,0,2,
/* out0493_em-eta13-phi24*/	9,6,0,3,6,1,3,6,2,4,61,1,1,61,2,1,62,0,2,62,1,3,67,0,1,67,2,2,
/* out0494_em-eta14-phi24*/	5,5,1,1,6,0,4,6,2,2,61,1,5,61,2,3,
/* out0495_em-eta15-phi24*/	5,1,0,1,5,1,2,5,2,4,61,0,4,61,1,3,
/* out0496_em-eta16-phi24*/	3,5,2,6,60,2,2,61,0,3,
/* out0497_em-eta17-phi24*/	4,0,1,4,5,2,2,60,0,6,60,2,3,
/* out0498_em-eta18-phi24*/	3,0,1,1,60,0,1,60,1,3,
/* out0499_em-eta19-phi24*/	0,
/* out0500_em-eta0-phi25*/	0,
/* out0501_em-eta1-phi25*/	0,
/* out0502_em-eta2-phi25*/	0,
/* out0503_em-eta3-phi25*/	0,
/* out0504_em-eta4-phi25*/	0,
/* out0505_em-eta5-phi25*/	0,
/* out0506_em-eta6-phi25*/	0,
/* out0507_em-eta7-phi25*/	0,
/* out0508_em-eta8-phi25*/	3,8,1,3,14,1,1,14,2,1,
/* out0509_em-eta9-phi25*/	8,8,0,4,8,1,10,8,2,6,63,2,1,64,0,12,64,2,3,69,1,5,69,2,1,
/* out0510_em-eta10-phi25*/	9,3,0,1,7,1,5,7,2,1,8,0,6,8,2,3,63,0,1,63,1,11,63,2,5,69,2,1,
/* out0511_em-eta11-phi25*/	7,7,0,1,7,1,2,7,2,11,62,1,1,62,2,3,63,0,7,63,1,3,
/* out0512_em-eta12-phi25*/	9,2,0,2,2,1,3,6,1,1,6,2,1,7,0,2,7,2,3,62,0,1,62,1,3,62,2,7,
/* out0513_em-eta13-phi25*/	3,2,0,3,6,2,7,62,0,10,
/* out0514_em-eta14-phi25*/	3,1,1,6,6,2,2,61,2,8,
/* out0515_em-eta15-phi25*/	4,1,0,6,1,1,1,61,0,4,61,2,3,
/* out0516_em-eta16-phi25*/	6,0,1,1,0,2,2,1,0,3,5,2,1,56,1,3,61,0,3,
/* out0517_em-eta17-phi25*/	4,0,1,5,0,2,2,56,1,3,60,0,5,
/* out0518_em-eta18-phi25*/	4,0,1,2,56,1,1,60,0,4,60,1,1,
/* out0519_em-eta19-phi25*/	0,
/* out0520_em-eta0-phi26*/	0,
/* out0521_em-eta1-phi26*/	0,
/* out0522_em-eta2-phi26*/	0,
/* out0523_em-eta3-phi26*/	0,
/* out0524_em-eta4-phi26*/	0,
/* out0525_em-eta5-phi26*/	0,
/* out0526_em-eta6-phi26*/	0,
/* out0527_em-eta7-phi26*/	0,
/* out0528_em-eta8-phi26*/	0,
/* out0529_em-eta9-phi26*/	7,3,1,1,4,0,12,4,2,3,8,2,6,59,1,3,64,0,4,64,2,13,
/* out0530_em-eta10-phi26*/	6,3,0,4,3,1,11,8,2,1,59,1,5,63,0,1,63,2,10,
/* out0531_em-eta11-phi26*/	6,2,1,3,3,0,9,7,2,1,58,1,7,62,2,1,63,0,7,
/* out0532_em-eta12-phi26*/	6,2,0,2,2,1,8,2,2,1,58,0,1,58,1,6,62,2,5,
/* out0533_em-eta13-phi26*/	5,2,0,9,2,2,1,57,1,6,57,2,1,62,0,3,
/* out0534_em-eta14-phi26*/	3,1,1,7,1,2,1,57,1,8,
/* out0535_em-eta15-phi26*/	9,1,0,2,1,1,1,1,2,3,56,1,1,56,2,2,57,0,2,57,1,1,61,0,1,61,2,1,
/* out0536_em-eta16-phi26*/	5,0,2,1,1,0,4,1,2,1,56,1,4,56,2,1,
/* out0537_em-eta17-phi26*/	3,0,2,6,56,0,1,56,1,4,
/* out0538_em-eta18-phi26*/	3,0,1,2,0,2,1,56,0,3,
/* out0539_em-eta19-phi26*/	0,
/* out0540_em-eta0-phi27*/	0,
/* out0541_em-eta1-phi27*/	0,
/* out0542_em-eta2-phi27*/	0,
/* out0543_em-eta3-phi27*/	0,
/* out0544_em-eta4-phi27*/	0,
/* out0545_em-eta5-phi27*/	0,
/* out0546_em-eta6-phi27*/	0,
/* out0547_em-eta7-phi27*/	0,
/* out0548_em-eta8-phi27*/	0,
/* out0549_em-eta9-phi27*/	5,3,1,1,4,0,4,4,2,13,59,1,4,59,2,11,
/* out0550_em-eta10-phi27*/	5,3,1,3,3,2,11,59,0,12,59,1,4,59,2,1,
/* out0551_em-eta11-phi27*/	5,2,1,1,3,0,2,3,2,5,58,1,2,58,2,12,
/* out0552_em-eta12-phi27*/	4,2,1,1,2,2,8,58,0,10,58,1,1,
/* out0553_em-eta13-phi27*/	3,2,2,6,57,2,9,58,0,1,
/* out0554_em-eta14-phi27*/	5,1,1,1,1,2,3,57,0,6,57,1,1,57,2,2,
/* out0555_em-eta15-phi27*/	3,1,2,6,56,2,3,57,0,4,
/* out0556_em-eta16-phi27*/	2,1,2,2,56,2,6,
/* out0557_em-eta17-phi27*/	3,0,2,2,56,0,4,56,2,1,
/* out0558_em-eta18-phi27*/	3,0,1,1,0,2,2,56,0,4,
/* out0559_em-eta19-phi27*/	0,
/* out0560_em-eta0-phi28*/	0,
/* out0561_em-eta1-phi28*/	0,
/* out0562_em-eta2-phi28*/	0,
/* out0563_em-eta3-phi28*/	0,
/* out0564_em-eta4-phi28*/	0,
/* out0565_em-eta5-phi28*/	0,
/* out0566_em-eta6-phi28*/	0,
/* out0567_em-eta7-phi28*/	0,
/* out0568_em-eta8-phi28*/	0,
/* out0569_em-eta9-phi28*/	1,59,2,3,
/* out0570_em-eta10-phi28*/	2,59,0,4,59,2,1,
/* out0571_em-eta11-phi28*/	1,58,2,4,
/* out0572_em-eta12-phi28*/	1,58,0,4,
/* out0573_em-eta13-phi28*/	1,57,2,2,
/* out0574_em-eta14-phi28*/	2,57,0,3,57,2,2,
/* out0575_em-eta15-phi28*/	1,57,0,1,
/* out0576_em-eta16-phi28*/	1,56,2,3,
/* out0577_em-eta17-phi28*/	1,56,0,3,
/* out0578_em-eta18-phi28*/	1,56,0,1,
/* out0579_em-eta19-phi28*/	0,
/* out0580_em-eta0-phi29*/	0,
/* out0581_em-eta1-phi29*/	0,
/* out0582_em-eta2-phi29*/	0,
/* out0583_em-eta3-phi29*/	0,
/* out0584_em-eta4-phi29*/	0,
/* out0585_em-eta5-phi29*/	0,
/* out0586_em-eta6-phi29*/	0,
/* out0587_em-eta7-phi29*/	0,
/* out0588_em-eta8-phi29*/	0,
/* out0589_em-eta9-phi29*/	0,
/* out0590_em-eta10-phi29*/	0,
/* out0591_em-eta11-phi29*/	0,
/* out0592_em-eta12-phi29*/	0,
/* out0593_em-eta13-phi29*/	0,
/* out0594_em-eta14-phi29*/	0,
/* out0595_em-eta15-phi29*/	0,
/* out0596_em-eta16-phi29*/	0,
/* out0597_em-eta17-phi29*/	0,
/* out0598_em-eta18-phi29*/	0,
/* out0599_em-eta19-phi29*/	0
};