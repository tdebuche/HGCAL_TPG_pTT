parameter integer matrixH [0:4356] = {
/* num inputs = 155(in0-in154) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 8 */
//* total number of input in adders 1292 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	1, 99, 0, 6, 
/* out0003_had-eta3-phi0*/	2, 98, 0, 3, 99, 0, 2, 
/* out0004_had-eta4-phi0*/	4, 87, 1, 1, 94, 0, 1, 94, 2, 5, 98, 0, 4, 
/* out0005_had-eta5-phi0*/	6, 86, 2, 1, 94, 0, 13, 94, 1, 11, 94, 2, 11, 97, 0, 4, 98, 0, 1, 
/* out0006_had-eta6-phi0*/	6, 86, 1, 1, 93, 0, 9, 93, 1, 3, 93, 2, 16, 94, 1, 5, 97, 0, 4, 
/* out0007_had-eta7-phi0*/	5, 92, 0, 2, 92, 2, 12, 93, 0, 2, 93, 1, 13, 96, 0, 3, 
/* out0008_had-eta8-phi0*/	4, 92, 0, 6, 92, 1, 9, 92, 2, 4, 96, 0, 3, 
/* out0009_had-eta9-phi0*/	4, 91, 0, 1, 91, 2, 11, 92, 1, 4, 96, 0, 2, 
/* out0010_had-eta10-phi0*/	4, 91, 0, 2, 91, 1, 9, 91, 2, 2, 95, 0, 6, 
/* out0011_had-eta11-phi0*/	3, 90, 2, 8, 91, 1, 3, 95, 0, 2, 
/* out0012_had-eta12-phi0*/	3, 90, 0, 1, 90, 1, 5, 90, 2, 4, 
/* out0013_had-eta13-phi0*/	2, 89, 2, 2, 90, 1, 6, 
/* out0014_had-eta14-phi0*/	1, 89, 2, 7, 
/* out0015_had-eta15-phi0*/	2, 89, 1, 4, 89, 2, 2, 
/* out0016_had-eta16-phi0*/	2, 88, 1, 1, 89, 1, 6, 
/* out0017_had-eta17-phi0*/	1, 88, 1, 4, 
/* out0018_had-eta18-phi0*/	1, 88, 1, 3, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	1, 99, 0, 6, 
/* out0023_had-eta3-phi1*/	2, 98, 0, 3, 99, 0, 2, 
/* out0024_had-eta4-phi1*/	3, 87, 0, 10, 87, 1, 6, 98, 0, 4, 
/* out0025_had-eta5-phi1*/	7, 86, 0, 5, 86, 2, 15, 87, 0, 3, 87, 1, 9, 94, 0, 2, 97, 0, 4, 98, 0, 1, 
/* out0026_had-eta6-phi1*/	5, 85, 2, 6, 86, 0, 2, 86, 1, 15, 93, 0, 4, 97, 0, 4, 
/* out0027_had-eta7-phi1*/	6, 85, 0, 1, 85, 1, 10, 85, 2, 9, 92, 0, 1, 93, 0, 1, 96, 0, 3, 
/* out0028_had-eta8-phi1*/	4, 84, 2, 9, 85, 1, 3, 92, 0, 7, 96, 0, 3, 
/* out0029_had-eta9-phi1*/	6, 84, 1, 8, 84, 2, 2, 91, 0, 5, 91, 2, 3, 92, 1, 3, 96, 0, 2, 
/* out0030_had-eta10-phi1*/	4, 83, 2, 5, 91, 0, 8, 91, 1, 3, 95, 0, 6, 
/* out0031_had-eta11-phi1*/	6, 83, 1, 3, 83, 2, 1, 90, 0, 4, 90, 2, 4, 91, 1, 1, 95, 0, 2, 
/* out0032_had-eta12-phi1*/	2, 90, 0, 8, 90, 1, 1, 
/* out0033_had-eta13-phi1*/	5, 82, 2, 1, 89, 0, 1, 89, 2, 2, 90, 0, 2, 90, 1, 4, 
/* out0034_had-eta14-phi1*/	2, 89, 0, 4, 89, 2, 2, 
/* out0035_had-eta15-phi1*/	3, 89, 0, 4, 89, 1, 1, 89, 2, 1, 
/* out0036_had-eta16-phi1*/	3, 88, 1, 1, 89, 0, 1, 89, 1, 4, 
/* out0037_had-eta17-phi1*/	2, 88, 0, 1, 88, 1, 4, 
/* out0038_had-eta18-phi1*/	2, 88, 0, 2, 88, 1, 2, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	1, 104, 0, 6, 
/* out0043_had-eta3-phi2*/	2, 103, 0, 3, 104, 0, 2, 
/* out0044_had-eta4-phi2*/	4, 80, 0, 2, 80, 2, 10, 87, 0, 3, 103, 0, 4, 
/* out0045_had-eta5-phi2*/	7, 79, 2, 4, 80, 0, 4, 80, 1, 15, 80, 2, 6, 86, 0, 5, 102, 0, 4, 103, 0, 1, 
/* out0046_had-eta6-phi2*/	6, 79, 1, 9, 79, 2, 9, 85, 0, 3, 85, 2, 1, 86, 0, 4, 102, 0, 4, 
/* out0047_had-eta7-phi2*/	5, 78, 2, 6, 79, 1, 1, 85, 0, 12, 85, 1, 2, 101, 0, 3, 
/* out0048_had-eta8-phi2*/	5, 78, 1, 3, 84, 0, 8, 84, 2, 5, 85, 1, 1, 101, 0, 3, 
/* out0049_had-eta9-phi2*/	4, 83, 2, 1, 84, 0, 6, 84, 1, 8, 101, 0, 2, 
/* out0050_had-eta10-phi2*/	3, 83, 0, 3, 83, 2, 9, 100, 0, 6, 
/* out0051_had-eta11-phi2*/	3, 83, 0, 1, 83, 1, 10, 100, 0, 2, 
/* out0052_had-eta12-phi2*/	3, 82, 2, 7, 83, 1, 1, 90, 0, 1, 
/* out0053_had-eta13-phi2*/	2, 82, 1, 4, 82, 2, 4, 
/* out0054_had-eta14-phi2*/	2, 82, 1, 4, 89, 0, 2, 
/* out0055_had-eta15-phi2*/	2, 81, 2, 2, 89, 0, 3, 
/* out0056_had-eta16-phi2*/	5, 81, 1, 1, 81, 2, 2, 88, 1, 1, 89, 0, 1, 89, 1, 1, 
/* out0057_had-eta17-phi2*/	2, 81, 1, 1, 88, 0, 6, 
/* out0058_had-eta18-phi2*/	1, 88, 0, 5, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	0, 
/* out0062_had-eta2-phi3*/	1, 104, 0, 6, 
/* out0063_had-eta3-phi3*/	2, 103, 0, 3, 104, 0, 2, 
/* out0064_had-eta4-phi3*/	3, 74, 2, 3, 80, 0, 2, 103, 0, 4, 
/* out0065_had-eta5-phi3*/	8, 74, 1, 9, 74, 2, 12, 79, 0, 3, 79, 2, 2, 80, 0, 8, 80, 1, 1, 102, 0, 4, 103, 0, 1, 
/* out0066_had-eta6-phi3*/	7, 73, 1, 1, 73, 2, 5, 74, 1, 1, 79, 0, 13, 79, 1, 5, 79, 2, 1, 102, 0, 4, 
/* out0067_had-eta7-phi3*/	6, 73, 1, 1, 78, 0, 9, 78, 1, 1, 78, 2, 10, 79, 1, 1, 101, 0, 3, 
/* out0068_had-eta8-phi3*/	5, 77, 2, 5, 78, 0, 1, 78, 1, 11, 84, 0, 1, 101, 0, 3, 
/* out0069_had-eta9-phi3*/	4, 77, 1, 5, 77, 2, 9, 84, 0, 1, 101, 0, 2, 
/* out0070_had-eta10-phi3*/	4, 76, 2, 1, 77, 1, 4, 83, 0, 7, 100, 0, 6, 
/* out0071_had-eta11-phi3*/	5, 76, 1, 1, 76, 2, 3, 83, 0, 5, 83, 1, 2, 100, 0, 2, 
/* out0072_had-eta12-phi3*/	2, 82, 0, 5, 82, 2, 3, 
/* out0073_had-eta13-phi3*/	3, 82, 0, 4, 82, 1, 3, 82, 2, 1, 
/* out0074_had-eta14-phi3*/	2, 81, 2, 2, 82, 1, 4, 
/* out0075_had-eta15-phi3*/	1, 81, 2, 5, 
/* out0076_had-eta16-phi3*/	2, 81, 1, 2, 81, 2, 2, 
/* out0077_had-eta17-phi3*/	1, 81, 1, 3, 
/* out0078_had-eta18-phi3*/	2, 81, 1, 1, 88, 0, 2, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	0, 
/* out0082_had-eta2-phi4*/	1, 109, 0, 6, 
/* out0083_had-eta3-phi4*/	2, 108, 0, 3, 109, 0, 2, 
/* out0084_had-eta4-phi4*/	3, 74, 0, 2, 74, 2, 1, 108, 0, 4, 
/* out0085_had-eta5-phi4*/	7, 73, 2, 1, 74, 0, 14, 74, 1, 5, 75, 1, 2, 75, 2, 8, 107, 0, 4, 108, 0, 1, 
/* out0086_had-eta6-phi4*/	6, 73, 0, 11, 73, 1, 5, 73, 2, 10, 74, 1, 1, 75, 1, 1, 107, 0, 4, 
/* out0087_had-eta7-phi4*/	4, 72, 2, 9, 73, 1, 9, 78, 0, 4, 106, 0, 3, 
/* out0088_had-eta8-phi4*/	7, 72, 1, 7, 72, 2, 4, 77, 0, 4, 77, 2, 1, 78, 0, 2, 78, 1, 1, 106, 0, 3, 
/* out0089_had-eta9-phi4*/	4, 77, 0, 12, 77, 1, 3, 77, 2, 1, 106, 0, 2, 
/* out0090_had-eta10-phi4*/	4, 76, 0, 1, 76, 2, 7, 77, 1, 4, 105, 0, 6, 
/* out0091_had-eta11-phi4*/	4, 76, 0, 1, 76, 1, 5, 76, 2, 5, 105, 0, 2, 
/* out0092_had-eta12-phi4*/	3, 60, 2, 1, 76, 1, 5, 82, 0, 3, 
/* out0093_had-eta13-phi4*/	2, 60, 2, 3, 82, 0, 4, 
/* out0094_had-eta14-phi4*/	5, 60, 1, 1, 60, 2, 1, 81, 0, 2, 81, 2, 1, 82, 1, 1, 
/* out0095_had-eta15-phi4*/	2, 81, 0, 4, 81, 2, 2, 
/* out0096_had-eta16-phi4*/	2, 81, 0, 2, 81, 1, 2, 
/* out0097_had-eta17-phi4*/	1, 81, 1, 4, 
/* out0098_had-eta18-phi4*/	0, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	0, 
/* out0102_had-eta2-phi5*/	1, 109, 0, 6, 
/* out0103_had-eta3-phi5*/	2, 108, 0, 3, 109, 0, 2, 
/* out0104_had-eta4-phi5*/	3, 75, 0, 1, 75, 2, 1, 108, 0, 4, 
/* out0105_had-eta5-phi5*/	5, 75, 0, 15, 75, 1, 8, 75, 2, 7, 107, 0, 4, 108, 0, 1, 
/* out0106_had-eta6-phi5*/	5, 68, 1, 1, 68, 2, 15, 73, 0, 4, 75, 1, 5, 107, 0, 4, 
/* out0107_had-eta7-phi5*/	6, 68, 1, 7, 68, 2, 1, 72, 0, 10, 72, 2, 3, 73, 0, 1, 106, 0, 3, 
/* out0108_had-eta8-phi5*/	4, 66, 2, 2, 72, 0, 6, 72, 1, 9, 106, 0, 3, 
/* out0109_had-eta9-phi5*/	3, 66, 1, 1, 66, 2, 13, 106, 0, 2, 
/* out0110_had-eta10-phi5*/	4, 66, 1, 6, 66, 2, 1, 76, 0, 6, 105, 0, 6, 
/* out0111_had-eta11-phi5*/	3, 76, 0, 8, 76, 1, 2, 105, 0, 2, 
/* out0112_had-eta12-phi5*/	2, 60, 2, 5, 76, 1, 3, 
/* out0113_had-eta13-phi5*/	2, 60, 1, 1, 60, 2, 6, 
/* out0114_had-eta14-phi5*/	1, 60, 1, 5, 
/* out0115_had-eta15-phi5*/	1, 81, 0, 4, 
/* out0116_had-eta16-phi5*/	1, 81, 0, 4, 
/* out0117_had-eta17-phi5*/	1, 81, 1, 2, 
/* out0118_had-eta18-phi5*/	0, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	0, 
/* out0122_had-eta2-phi6*/	1, 114, 0, 6, 
/* out0123_had-eta3-phi6*/	2, 113, 0, 3, 114, 0, 2, 
/* out0124_had-eta4-phi6*/	3, 70, 0, 1, 70, 2, 1, 113, 0, 4, 
/* out0125_had-eta5-phi6*/	5, 70, 0, 7, 70, 1, 8, 70, 2, 15, 112, 0, 4, 113, 0, 1, 
/* out0126_had-eta6-phi6*/	5, 68, 0, 15, 68, 1, 1, 69, 2, 4, 70, 1, 5, 112, 0, 4, 
/* out0127_had-eta7-phi6*/	6, 67, 0, 3, 67, 2, 10, 68, 0, 1, 68, 1, 7, 69, 2, 1, 111, 0, 3, 
/* out0128_had-eta8-phi6*/	4, 66, 0, 3, 67, 1, 9, 67, 2, 6, 111, 0, 3, 
/* out0129_had-eta9-phi6*/	3, 66, 0, 13, 66, 1, 2, 111, 0, 2, 
/* out0130_had-eta10-phi6*/	3, 61, 2, 6, 66, 1, 7, 110, 0, 6, 
/* out0131_had-eta11-phi6*/	3, 61, 1, 2, 61, 2, 8, 110, 0, 2, 
/* out0132_had-eta12-phi6*/	2, 60, 0, 5, 61, 1, 3, 
/* out0133_had-eta13-phi6*/	2, 60, 0, 6, 60, 1, 1, 
/* out0134_had-eta14-phi6*/	1, 60, 1, 6, 
/* out0135_had-eta15-phi6*/	2, 53, 2, 4, 60, 1, 1, 
/* out0136_had-eta16-phi6*/	1, 53, 2, 4, 
/* out0137_had-eta17-phi6*/	1, 53, 1, 2, 
/* out0138_had-eta18-phi6*/	0, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	0, 
/* out0142_had-eta2-phi7*/	1, 114, 0, 6, 
/* out0143_had-eta3-phi7*/	2, 113, 0, 3, 114, 0, 2, 
/* out0144_had-eta4-phi7*/	3, 71, 0, 1, 71, 2, 2, 113, 0, 4, 
/* out0145_had-eta5-phi7*/	7, 69, 0, 1, 70, 0, 8, 70, 1, 2, 71, 1, 5, 71, 2, 14, 112, 0, 4, 113, 0, 1, 
/* out0146_had-eta6-phi7*/	6, 69, 0, 10, 69, 1, 5, 69, 2, 11, 70, 1, 1, 71, 1, 1, 112, 0, 4, 
/* out0147_had-eta7-phi7*/	4, 63, 2, 4, 67, 0, 9, 69, 1, 9, 111, 0, 3, 
/* out0148_had-eta8-phi7*/	7, 62, 0, 1, 62, 2, 4, 63, 1, 1, 63, 2, 2, 67, 0, 4, 67, 1, 7, 111, 0, 3, 
/* out0149_had-eta9-phi7*/	4, 62, 0, 1, 62, 1, 3, 62, 2, 12, 111, 0, 2, 
/* out0150_had-eta10-phi7*/	4, 61, 0, 7, 61, 2, 1, 62, 1, 4, 110, 0, 6, 
/* out0151_had-eta11-phi7*/	4, 61, 0, 5, 61, 1, 5, 61, 2, 1, 110, 0, 2, 
/* out0152_had-eta12-phi7*/	3, 54, 2, 3, 60, 0, 1, 61, 1, 5, 
/* out0153_had-eta13-phi7*/	2, 54, 2, 4, 60, 0, 3, 
/* out0154_had-eta14-phi7*/	5, 53, 0, 1, 53, 2, 2, 54, 1, 1, 60, 0, 1, 60, 1, 1, 
/* out0155_had-eta15-phi7*/	2, 53, 0, 2, 53, 2, 4, 
/* out0156_had-eta16-phi7*/	2, 53, 1, 2, 53, 2, 2, 
/* out0157_had-eta17-phi7*/	1, 53, 1, 4, 
/* out0158_had-eta18-phi7*/	0, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	0, 
/* out0162_had-eta2-phi8*/	1, 119, 0, 6, 
/* out0163_had-eta3-phi8*/	2, 118, 0, 3, 119, 0, 2, 
/* out0164_had-eta4-phi8*/	3, 65, 2, 2, 71, 0, 3, 118, 0, 4, 
/* out0165_had-eta5-phi8*/	8, 64, 0, 2, 64, 2, 3, 65, 1, 1, 65, 2, 8, 71, 0, 12, 71, 1, 9, 117, 0, 4, 118, 0, 1, 
/* out0166_had-eta6-phi8*/	7, 64, 0, 1, 64, 1, 5, 64, 2, 13, 69, 0, 5, 69, 1, 1, 71, 1, 1, 117, 0, 4, 
/* out0167_had-eta7-phi8*/	6, 63, 0, 10, 63, 1, 1, 63, 2, 9, 64, 1, 1, 69, 1, 1, 116, 0, 3, 
/* out0168_had-eta8-phi8*/	5, 56, 2, 1, 62, 0, 5, 63, 1, 11, 63, 2, 1, 116, 0, 3, 
/* out0169_had-eta9-phi8*/	4, 56, 2, 1, 62, 0, 9, 62, 1, 5, 116, 0, 2, 
/* out0170_had-eta10-phi8*/	4, 55, 2, 7, 61, 0, 1, 62, 1, 4, 115, 0, 6, 
/* out0171_had-eta11-phi8*/	5, 55, 1, 2, 55, 2, 5, 61, 0, 3, 61, 1, 1, 115, 0, 2, 
/* out0172_had-eta12-phi8*/	2, 54, 0, 3, 54, 2, 5, 
/* out0173_had-eta13-phi8*/	3, 54, 0, 1, 54, 1, 3, 54, 2, 4, 
/* out0174_had-eta14-phi8*/	2, 53, 0, 2, 54, 1, 4, 
/* out0175_had-eta15-phi8*/	1, 53, 0, 5, 
/* out0176_had-eta16-phi8*/	2, 53, 0, 2, 53, 1, 2, 
/* out0177_had-eta17-phi8*/	1, 53, 1, 3, 
/* out0178_had-eta18-phi8*/	2, 46, 1, 2, 53, 1, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	0, 
/* out0182_had-eta2-phi9*/	1, 119, 0, 6, 
/* out0183_had-eta3-phi9*/	2, 118, 0, 3, 119, 0, 2, 
/* out0184_had-eta4-phi9*/	4, 59, 1, 3, 65, 0, 10, 65, 2, 2, 118, 0, 4, 
/* out0185_had-eta5-phi9*/	7, 58, 2, 5, 64, 0, 4, 65, 0, 6, 65, 1, 15, 65, 2, 4, 117, 0, 4, 118, 0, 1, 
/* out0186_had-eta6-phi9*/	6, 57, 0, 1, 57, 2, 3, 58, 2, 4, 64, 0, 9, 64, 1, 9, 117, 0, 4, 
/* out0187_had-eta7-phi9*/	5, 57, 1, 2, 57, 2, 12, 63, 0, 6, 64, 1, 1, 116, 0, 3, 
/* out0188_had-eta8-phi9*/	5, 56, 0, 5, 56, 2, 8, 57, 1, 1, 63, 1, 3, 116, 0, 3, 
/* out0189_had-eta9-phi9*/	4, 55, 0, 1, 56, 1, 8, 56, 2, 6, 116, 0, 2, 
/* out0190_had-eta10-phi9*/	3, 55, 0, 9, 55, 2, 3, 115, 0, 6, 
/* out0191_had-eta11-phi9*/	3, 55, 1, 10, 55, 2, 1, 115, 0, 2, 
/* out0192_had-eta12-phi9*/	3, 48, 2, 1, 54, 0, 7, 55, 1, 1, 
/* out0193_had-eta13-phi9*/	2, 54, 0, 4, 54, 1, 4, 
/* out0194_had-eta14-phi9*/	2, 47, 2, 2, 54, 1, 4, 
/* out0195_had-eta15-phi9*/	2, 47, 2, 3, 53, 0, 2, 
/* out0196_had-eta16-phi9*/	3, 47, 2, 1, 53, 0, 2, 53, 1, 1, 
/* out0197_had-eta17-phi9*/	2, 46, 1, 6, 53, 1, 1, 
/* out0198_had-eta18-phi9*/	1, 46, 1, 5, 
/* out0199_had-eta19-phi9*/	0, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	0, 
/* out0202_had-eta2-phi10*/	1, 124, 0, 6, 
/* out0203_had-eta3-phi10*/	2, 123, 0, 3, 124, 0, 2, 
/* out0204_had-eta4-phi10*/	3, 59, 0, 6, 59, 1, 10, 123, 0, 4, 
/* out0205_had-eta5-phi10*/	7, 52, 2, 2, 58, 0, 15, 58, 2, 5, 59, 0, 9, 59, 1, 3, 122, 0, 4, 123, 0, 1, 
/* out0206_had-eta6-phi10*/	5, 51, 2, 4, 57, 0, 6, 58, 1, 15, 58, 2, 2, 122, 0, 4, 
/* out0207_had-eta7-phi10*/	6, 50, 2, 1, 51, 2, 1, 57, 0, 9, 57, 1, 10, 57, 2, 1, 121, 0, 3, 
/* out0208_had-eta8-phi10*/	4, 50, 2, 7, 56, 0, 9, 57, 1, 3, 121, 0, 3, 
/* out0209_had-eta9-phi10*/	4, 49, 2, 5, 56, 0, 2, 56, 1, 8, 121, 0, 2, 
/* out0210_had-eta10-phi10*/	3, 49, 2, 8, 55, 0, 5, 120, 0, 6, 
/* out0211_had-eta11-phi10*/	5, 48, 0, 1, 48, 2, 4, 55, 0, 1, 55, 1, 3, 120, 0, 2, 
/* out0212_had-eta12-phi10*/	1, 48, 2, 8, 
/* out0213_had-eta13-phi10*/	5, 47, 0, 1, 47, 2, 1, 48, 1, 2, 48, 2, 2, 54, 0, 1, 
/* out0214_had-eta14-phi10*/	2, 47, 0, 2, 47, 2, 4, 
/* out0215_had-eta15-phi10*/	2, 47, 1, 1, 47, 2, 4, 
/* out0216_had-eta16-phi10*/	3, 46, 0, 1, 47, 1, 3, 47, 2, 1, 
/* out0217_had-eta17-phi10*/	2, 46, 0, 3, 46, 1, 1, 
/* out0218_had-eta18-phi10*/	2, 46, 0, 1, 46, 1, 2, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	0, 
/* out0222_had-eta2-phi11*/	1, 124, 0, 6, 
/* out0223_had-eta3-phi11*/	2, 123, 0, 3, 124, 0, 2, 
/* out0224_had-eta4-phi11*/	4, 52, 0, 5, 52, 2, 1, 59, 0, 1, 123, 0, 4, 
/* out0225_had-eta5-phi11*/	6, 52, 0, 7, 52, 1, 11, 52, 2, 13, 58, 0, 1, 122, 0, 4, 123, 0, 1, 
/* out0226_had-eta6-phi11*/	6, 51, 0, 12, 51, 1, 3, 51, 2, 9, 52, 1, 1, 58, 1, 1, 122, 0, 4, 
/* out0227_had-eta7-phi11*/	5, 50, 0, 8, 50, 2, 2, 51, 1, 9, 51, 2, 2, 121, 0, 3, 
/* out0228_had-eta8-phi11*/	4, 50, 0, 4, 50, 1, 9, 50, 2, 6, 121, 0, 3, 
/* out0229_had-eta9-phi11*/	4, 49, 0, 10, 49, 2, 1, 50, 1, 3, 121, 0, 2, 
/* out0230_had-eta10-phi11*/	4, 49, 0, 2, 49, 1, 9, 49, 2, 2, 120, 0, 6, 
/* out0231_had-eta11-phi11*/	3, 48, 0, 8, 49, 1, 3, 120, 0, 2, 
/* out0232_had-eta12-phi11*/	3, 48, 0, 3, 48, 1, 5, 48, 2, 1, 
/* out0233_had-eta13-phi11*/	2, 47, 0, 2, 48, 1, 5, 
/* out0234_had-eta14-phi11*/	1, 47, 0, 6, 
/* out0235_had-eta15-phi11*/	2, 47, 0, 1, 47, 1, 4, 
/* out0236_had-eta16-phi11*/	1, 47, 1, 4, 
/* out0237_had-eta17-phi11*/	1, 46, 0, 4, 
/* out0238_had-eta18-phi11*/	1, 46, 0, 3, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	0, 
/* out0242_had-eta2-phi12*/	1, 129, 0, 6, 
/* out0243_had-eta3-phi12*/	2, 128, 0, 3, 129, 0, 2, 
/* out0244_had-eta4-phi12*/	3, 45, 0, 3, 45, 1, 9, 128, 0, 4, 
/* out0245_had-eta5-phi12*/	8, 44, 0, 8, 44, 2, 7, 45, 0, 6, 45, 1, 7, 52, 0, 4, 52, 1, 4, 127, 0, 4, 128, 0, 1, 
/* out0246_had-eta6-phi12*/	7, 43, 0, 3, 43, 2, 1, 44, 1, 7, 44, 2, 9, 51, 0, 4, 51, 1, 2, 127, 0, 4, 
/* out0247_had-eta7-phi12*/	6, 43, 0, 3, 43, 1, 2, 43, 2, 14, 50, 0, 1, 51, 1, 2, 126, 0, 3, 
/* out0248_had-eta8-phi12*/	7, 42, 0, 3, 42, 2, 5, 43, 1, 2, 43, 2, 1, 50, 0, 3, 50, 1, 4, 126, 0, 3, 
/* out0249_had-eta9-phi12*/	4, 42, 1, 1, 42, 2, 11, 49, 0, 3, 126, 0, 2, 
/* out0250_had-eta10-phi12*/	6, 41, 0, 1, 41, 2, 5, 42, 1, 1, 49, 0, 1, 49, 1, 4, 125, 0, 6, 
/* out0251_had-eta11-phi12*/	3, 41, 2, 8, 48, 0, 2, 125, 0, 2, 
/* out0252_had-eta12-phi12*/	5, 40, 2, 2, 41, 1, 1, 41, 2, 1, 48, 0, 2, 48, 1, 3, 
/* out0253_had-eta13-phi12*/	2, 40, 2, 6, 48, 1, 1, 
/* out0254_had-eta14-phi12*/	2, 40, 2, 3, 47, 0, 3, 
/* out0255_had-eta15-phi12*/	3, 39, 2, 1, 47, 0, 1, 47, 1, 3, 
/* out0256_had-eta16-phi12*/	2, 39, 2, 3, 47, 1, 1, 
/* out0257_had-eta17-phi12*/	2, 39, 2, 3, 46, 0, 1, 
/* out0258_had-eta18-phi12*/	1, 46, 0, 3, 
/* out0259_had-eta19-phi12*/	0, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	0, 
/* out0262_had-eta2-phi13*/	1, 129, 0, 6, 
/* out0263_had-eta3-phi13*/	2, 128, 0, 3, 129, 0, 2, 
/* out0264_had-eta4-phi13*/	4, 38, 0, 5, 38, 2, 2, 45, 0, 4, 128, 0, 4, 
/* out0265_had-eta5-phi13*/	8, 37, 0, 1, 38, 0, 2, 38, 1, 4, 38, 2, 14, 44, 0, 8, 45, 0, 3, 127, 0, 4, 128, 0, 1, 
/* out0266_had-eta6-phi13*/	5, 37, 0, 2, 37, 2, 12, 43, 0, 3, 44, 1, 9, 127, 0, 4, 
/* out0267_had-eta7-phi13*/	6, 36, 2, 3, 37, 1, 1, 37, 2, 2, 43, 0, 7, 43, 1, 9, 126, 0, 3, 
/* out0268_had-eta8-phi13*/	4, 36, 2, 5, 42, 0, 11, 43, 1, 3, 126, 0, 3, 
/* out0269_had-eta9-phi13*/	4, 35, 2, 1, 42, 0, 2, 42, 1, 12, 126, 0, 2, 
/* out0270_had-eta10-phi13*/	3, 41, 0, 11, 42, 1, 1, 125, 0, 6, 
/* out0271_had-eta11-phi13*/	4, 41, 0, 1, 41, 1, 8, 41, 2, 2, 125, 0, 2, 
/* out0272_had-eta12-phi13*/	2, 40, 0, 6, 41, 1, 3, 
/* out0273_had-eta13-phi13*/	3, 40, 0, 3, 40, 1, 1, 40, 2, 3, 
/* out0274_had-eta14-phi13*/	2, 40, 1, 4, 40, 2, 2, 
/* out0275_had-eta15-phi13*/	3, 39, 0, 3, 39, 2, 1, 40, 1, 1, 
/* out0276_had-eta16-phi13*/	2, 39, 0, 1, 39, 2, 4, 
/* out0277_had-eta17-phi13*/	1, 39, 2, 3, 
/* out0278_had-eta18-phi13*/	2, 39, 1, 1, 39, 2, 1, 
/* out0279_had-eta19-phi13*/	0, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	0, 
/* out0282_had-eta2-phi14*/	1, 134, 0, 6, 
/* out0283_had-eta3-phi14*/	2, 133, 0, 3, 134, 0, 2, 
/* out0284_had-eta4-phi14*/	2, 38, 0, 5, 133, 0, 4, 
/* out0285_had-eta5-phi14*/	7, 32, 0, 2, 32, 2, 11, 37, 0, 2, 38, 0, 4, 38, 1, 12, 132, 0, 4, 133, 0, 1, 
/* out0286_had-eta6-phi14*/	6, 31, 2, 1, 32, 2, 2, 37, 0, 11, 37, 1, 10, 37, 2, 2, 132, 0, 4, 
/* out0287_had-eta7-phi14*/	5, 31, 2, 2, 36, 0, 13, 36, 2, 2, 37, 1, 5, 131, 0, 3, 
/* out0288_had-eta8-phi14*/	4, 35, 0, 1, 36, 1, 10, 36, 2, 6, 131, 0, 3, 
/* out0289_had-eta9-phi14*/	4, 35, 0, 6, 35, 2, 8, 42, 1, 1, 131, 0, 2, 
/* out0290_had-eta10-phi14*/	4, 35, 1, 3, 35, 2, 7, 41, 0, 3, 130, 0, 6, 
/* out0291_had-eta11-phi14*/	4, 34, 0, 1, 34, 2, 5, 41, 1, 4, 130, 0, 2, 
/* out0292_had-eta12-phi14*/	2, 34, 2, 5, 40, 0, 3, 
/* out0293_had-eta13-phi14*/	2, 40, 0, 4, 40, 1, 4, 
/* out0294_had-eta14-phi14*/	2, 33, 2, 1, 40, 1, 5, 
/* out0295_had-eta15-phi14*/	1, 39, 0, 5, 
/* out0296_had-eta16-phi14*/	2, 39, 0, 3, 39, 1, 1, 
/* out0297_had-eta17-phi14*/	1, 39, 1, 4, 
/* out0298_had-eta18-phi14*/	1, 39, 1, 2, 
/* out0299_had-eta19-phi14*/	0, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	0, 
/* out0302_had-eta2-phi15*/	1, 134, 0, 6, 
/* out0303_had-eta3-phi15*/	2, 133, 0, 3, 134, 0, 2, 
/* out0304_had-eta4-phi15*/	2, 28, 1, 10, 133, 0, 4, 
/* out0305_had-eta5-phi15*/	7, 26, 2, 2, 28, 1, 5, 32, 0, 14, 32, 1, 10, 32, 2, 2, 132, 0, 4, 133, 0, 1, 
/* out0306_had-eta6-phi15*/	7, 26, 2, 1, 31, 0, 13, 31, 1, 1, 31, 2, 5, 32, 1, 6, 32, 2, 1, 132, 0, 4, 
/* out0307_had-eta7-phi15*/	6, 30, 0, 3, 31, 1, 7, 31, 2, 8, 36, 0, 3, 36, 1, 1, 131, 0, 3, 
/* out0308_had-eta8-phi15*/	5, 30, 0, 1, 30, 2, 11, 35, 0, 1, 36, 1, 5, 131, 0, 3, 
/* out0309_had-eta9-phi15*/	4, 30, 2, 2, 35, 0, 8, 35, 1, 5, 131, 0, 2, 
/* out0310_had-eta10-phi15*/	4, 29, 2, 1, 34, 0, 3, 35, 1, 8, 130, 0, 6, 
/* out0311_had-eta11-phi15*/	4, 34, 0, 8, 34, 1, 1, 34, 2, 2, 130, 0, 2, 
/* out0312_had-eta12-phi15*/	2, 34, 1, 5, 34, 2, 4, 
/* out0313_had-eta13-phi15*/	4, 33, 0, 3, 33, 2, 2, 34, 1, 1, 40, 1, 1, 
/* out0314_had-eta14-phi15*/	1, 33, 2, 6, 
/* out0315_had-eta15-phi15*/	2, 33, 2, 3, 39, 0, 2, 
/* out0316_had-eta16-phi15*/	2, 39, 0, 2, 39, 1, 2, 
/* out0317_had-eta17-phi15*/	1, 39, 1, 4, 
/* out0318_had-eta18-phi15*/	1, 39, 1, 1, 
/* out0319_had-eta19-phi15*/	0, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	0, 
/* out0322_had-eta2-phi16*/	1, 139, 0, 6, 
/* out0323_had-eta3-phi16*/	2, 138, 0, 3, 139, 0, 2, 
/* out0324_had-eta4-phi16*/	4, 27, 1, 3, 28, 0, 8, 28, 1, 1, 138, 0, 4, 
/* out0325_had-eta5-phi16*/	7, 26, 0, 14, 26, 1, 3, 26, 2, 6, 27, 1, 4, 28, 0, 8, 137, 0, 4, 138, 0, 1, 
/* out0326_had-eta6-phi16*/	7, 25, 0, 4, 25, 2, 2, 26, 1, 7, 26, 2, 7, 31, 0, 3, 31, 1, 3, 137, 0, 4, 
/* out0327_had-eta7-phi16*/	4, 25, 2, 11, 30, 0, 6, 31, 1, 5, 136, 0, 3, 
/* out0328_had-eta8-phi16*/	4, 30, 0, 6, 30, 1, 10, 30, 2, 2, 136, 0, 3, 
/* out0329_had-eta9-phi16*/	5, 29, 0, 8, 29, 2, 3, 30, 1, 4, 30, 2, 1, 136, 0, 2, 
/* out0330_had-eta10-phi16*/	3, 29, 1, 1, 29, 2, 11, 135, 0, 6, 
/* out0331_had-eta11-phi16*/	6, 14, 2, 1, 29, 1, 1, 29, 2, 1, 34, 0, 4, 34, 1, 3, 135, 0, 2, 
/* out0332_had-eta12-phi16*/	3, 14, 2, 2, 33, 0, 1, 34, 1, 6, 
/* out0333_had-eta13-phi16*/	1, 33, 0, 7, 
/* out0334_had-eta14-phi16*/	3, 33, 0, 1, 33, 1, 3, 33, 2, 2, 
/* out0335_had-eta15-phi16*/	2, 33, 1, 3, 33, 2, 2, 
/* out0336_had-eta16-phi16*/	3, 0, 0, 1, 0, 2, 2, 39, 1, 1, 
/* out0337_had-eta17-phi16*/	1, 0, 2, 5, 
/* out0338_had-eta18-phi16*/	1, 0, 2, 2, 
/* out0339_had-eta19-phi16*/	0, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	0, 
/* out0342_had-eta2-phi17*/	1, 139, 0, 6, 
/* out0343_had-eta3-phi17*/	2, 138, 0, 3, 139, 0, 2, 
/* out0344_had-eta4-phi17*/	3, 27, 0, 4, 27, 1, 2, 138, 0, 4, 
/* out0345_had-eta5-phi17*/	8, 23, 0, 8, 23, 2, 5, 26, 0, 2, 26, 1, 3, 27, 0, 12, 27, 1, 7, 137, 0, 4, 138, 0, 1, 
/* out0346_had-eta6-phi17*/	5, 23, 2, 11, 25, 0, 11, 25, 1, 1, 26, 1, 3, 137, 0, 4, 
/* out0347_had-eta7-phi17*/	5, 19, 0, 2, 25, 0, 1, 25, 1, 15, 25, 2, 3, 136, 0, 3, 
/* out0348_had-eta8-phi17*/	4, 19, 0, 5, 19, 2, 10, 30, 1, 2, 136, 0, 3, 
/* out0349_had-eta9-phi17*/	4, 19, 2, 6, 29, 0, 8, 29, 1, 2, 136, 0, 2, 
/* out0350_had-eta10-phi17*/	2, 29, 1, 11, 135, 0, 6, 
/* out0351_had-eta11-phi17*/	4, 14, 0, 7, 14, 2, 2, 29, 1, 1, 135, 0, 2, 
/* out0352_had-eta12-phi17*/	1, 14, 2, 9, 
/* out0353_had-eta13-phi17*/	3, 14, 2, 2, 33, 0, 4, 33, 1, 1, 
/* out0354_had-eta14-phi17*/	1, 33, 1, 6, 
/* out0355_had-eta15-phi17*/	2, 0, 0, 2, 33, 1, 3, 
/* out0356_had-eta16-phi17*/	1, 0, 0, 4, 
/* out0357_had-eta17-phi17*/	1, 0, 2, 4, 
/* out0358_had-eta18-phi17*/	1, 0, 2, 3, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	0, 
/* out0362_had-eta2-phi18*/	1, 144, 0, 6, 
/* out0363_had-eta3-phi18*/	2, 143, 0, 3, 144, 0, 2, 
/* out0364_had-eta4-phi18*/	3, 24, 0, 2, 24, 1, 4, 143, 0, 4, 
/* out0365_had-eta5-phi18*/	8, 21, 0, 2, 21, 2, 3, 23, 0, 8, 23, 1, 5, 24, 0, 7, 24, 1, 12, 142, 0, 4, 143, 0, 1, 
/* out0366_had-eta6-phi18*/	5, 20, 0, 11, 20, 2, 1, 21, 2, 3, 23, 1, 11, 142, 0, 4, 
/* out0367_had-eta7-phi18*/	5, 19, 0, 3, 20, 0, 1, 20, 1, 3, 20, 2, 15, 141, 0, 3, 
/* out0368_had-eta8-phi18*/	4, 16, 2, 2, 19, 0, 6, 19, 1, 10, 141, 0, 3, 
/* out0369_had-eta9-phi18*/	4, 15, 0, 8, 15, 2, 2, 19, 1, 6, 141, 0, 2, 
/* out0370_had-eta10-phi18*/	3, 14, 0, 1, 15, 2, 11, 140, 0, 6, 
/* out0371_had-eta11-phi18*/	4, 14, 0, 8, 14, 1, 2, 15, 2, 1, 140, 0, 2, 
/* out0372_had-eta12-phi18*/	1, 14, 1, 8, 
/* out0373_had-eta13-phi18*/	3, 1, 0, 4, 1, 2, 1, 14, 1, 3, 
/* out0374_had-eta14-phi18*/	1, 1, 2, 6, 
/* out0375_had-eta15-phi18*/	2, 0, 0, 2, 1, 2, 3, 
/* out0376_had-eta16-phi18*/	1, 0, 0, 4, 
/* out0377_had-eta17-phi18*/	2, 0, 0, 1, 0, 1, 4, 
/* out0378_had-eta18-phi18*/	1, 0, 1, 2, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	0, 
/* out0382_had-eta2-phi19*/	1, 144, 0, 6, 
/* out0383_had-eta3-phi19*/	2, 143, 0, 3, 144, 0, 2, 
/* out0384_had-eta4-phi19*/	4, 22, 0, 1, 22, 1, 8, 24, 0, 3, 143, 0, 4, 
/* out0385_had-eta5-phi19*/	7, 21, 0, 14, 21, 1, 6, 21, 2, 3, 22, 1, 8, 24, 0, 4, 142, 0, 4, 143, 0, 1, 
/* out0386_had-eta6-phi19*/	7, 17, 0, 3, 17, 2, 3, 20, 0, 4, 20, 1, 2, 21, 1, 7, 21, 2, 7, 142, 0, 4, 
/* out0387_had-eta7-phi19*/	4, 16, 0, 6, 17, 2, 5, 20, 1, 11, 141, 0, 3, 
/* out0388_had-eta8-phi19*/	4, 16, 0, 6, 16, 1, 2, 16, 2, 10, 141, 0, 3, 
/* out0389_had-eta9-phi19*/	5, 15, 0, 8, 15, 1, 3, 16, 1, 1, 16, 2, 4, 141, 0, 2, 
/* out0390_had-eta10-phi19*/	3, 15, 1, 11, 15, 2, 1, 140, 0, 6, 
/* out0391_had-eta11-phi19*/	6, 2, 0, 4, 2, 2, 3, 14, 1, 1, 15, 1, 1, 15, 2, 1, 140, 0, 2, 
/* out0392_had-eta12-phi19*/	3, 1, 0, 1, 2, 2, 6, 14, 1, 2, 
/* out0393_had-eta13-phi19*/	1, 1, 0, 7, 
/* out0394_had-eta14-phi19*/	3, 1, 0, 1, 1, 1, 2, 1, 2, 3, 
/* out0395_had-eta15-phi19*/	2, 1, 1, 2, 1, 2, 3, 
/* out0396_had-eta16-phi19*/	3, 0, 0, 2, 0, 1, 3, 7, 2, 1, 
/* out0397_had-eta17-phi19*/	1, 0, 1, 5, 
/* out0398_had-eta18-phi19*/	1, 0, 1, 2, 
/* out0399_had-eta19-phi19*/	0, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	0, 
/* out0402_had-eta2-phi20*/	1, 149, 0, 6, 
/* out0403_had-eta3-phi20*/	2, 148, 0, 3, 149, 0, 2, 
/* out0404_had-eta4-phi20*/	2, 22, 0, 10, 148, 0, 4, 
/* out0405_had-eta5-phi20*/	7, 18, 0, 14, 18, 1, 2, 18, 2, 10, 21, 1, 2, 22, 0, 5, 147, 0, 4, 148, 0, 1, 
/* out0406_had-eta6-phi20*/	7, 17, 0, 13, 17, 1, 5, 17, 2, 1, 18, 1, 1, 18, 2, 6, 21, 1, 1, 147, 0, 4, 
/* out0407_had-eta7-phi20*/	6, 4, 0, 3, 4, 2, 1, 16, 0, 3, 17, 1, 8, 17, 2, 7, 146, 0, 3, 
/* out0408_had-eta8-phi20*/	5, 3, 0, 1, 4, 2, 5, 16, 0, 1, 16, 1, 11, 146, 0, 3, 
/* out0409_had-eta9-phi20*/	4, 3, 0, 8, 3, 2, 5, 16, 1, 2, 146, 0, 2, 
/* out0410_had-eta10-phi20*/	4, 2, 0, 3, 3, 2, 8, 15, 1, 1, 145, 0, 6, 
/* out0411_had-eta11-phi20*/	4, 2, 0, 8, 2, 1, 2, 2, 2, 1, 145, 0, 2, 
/* out0412_had-eta12-phi20*/	2, 2, 1, 4, 2, 2, 5, 
/* out0413_had-eta13-phi20*/	4, 1, 0, 3, 1, 1, 2, 2, 2, 1, 8, 2, 1, 
/* out0414_had-eta14-phi20*/	1, 1, 1, 6, 
/* out0415_had-eta15-phi20*/	2, 1, 1, 3, 7, 0, 2, 
/* out0416_had-eta16-phi20*/	2, 7, 0, 2, 7, 2, 2, 
/* out0417_had-eta17-phi20*/	1, 7, 2, 4, 
/* out0418_had-eta18-phi20*/	1, 7, 2, 1, 
/* out0419_had-eta19-phi20*/	0, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	0, 
/* out0422_had-eta2-phi21*/	1, 149, 0, 6, 
/* out0423_had-eta3-phi21*/	2, 148, 0, 3, 149, 0, 2, 
/* out0424_had-eta4-phi21*/	2, 6, 0, 5, 148, 0, 4, 
/* out0425_had-eta5-phi21*/	7, 5, 0, 2, 6, 0, 4, 6, 2, 12, 18, 0, 2, 18, 1, 11, 147, 0, 4, 148, 0, 1, 
/* out0426_had-eta6-phi21*/	6, 5, 0, 11, 5, 1, 2, 5, 2, 10, 17, 1, 1, 18, 1, 2, 147, 0, 4, 
/* out0427_had-eta7-phi21*/	5, 4, 0, 13, 4, 1, 2, 5, 2, 5, 17, 1, 2, 146, 0, 3, 
/* out0428_had-eta8-phi21*/	4, 3, 0, 1, 4, 1, 6, 4, 2, 10, 146, 0, 3, 
/* out0429_had-eta9-phi21*/	4, 3, 0, 6, 3, 1, 8, 10, 2, 1, 146, 0, 2, 
/* out0430_had-eta10-phi21*/	4, 3, 1, 7, 3, 2, 3, 9, 0, 3, 145, 0, 6, 
/* out0431_had-eta11-phi21*/	4, 2, 0, 1, 2, 1, 5, 9, 2, 4, 145, 0, 2, 
/* out0432_had-eta12-phi21*/	2, 2, 1, 5, 8, 0, 3, 
/* out0433_had-eta13-phi21*/	2, 8, 0, 4, 8, 2, 4, 
/* out0434_had-eta14-phi21*/	2, 1, 1, 1, 8, 2, 5, 
/* out0435_had-eta15-phi21*/	1, 7, 0, 5, 
/* out0436_had-eta16-phi21*/	2, 7, 0, 3, 7, 2, 1, 
/* out0437_had-eta17-phi21*/	1, 7, 2, 4, 
/* out0438_had-eta18-phi21*/	1, 7, 2, 2, 
/* out0439_had-eta19-phi21*/	0, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	0, 
/* out0442_had-eta2-phi22*/	1, 154, 0, 6, 
/* out0443_had-eta3-phi22*/	2, 153, 0, 3, 154, 0, 2, 
/* out0444_had-eta4-phi22*/	4, 6, 0, 5, 6, 1, 2, 13, 1, 4, 153, 0, 4, 
/* out0445_had-eta5-phi22*/	8, 5, 0, 1, 6, 0, 2, 6, 1, 14, 6, 2, 4, 12, 0, 8, 13, 1, 3, 152, 0, 4, 153, 0, 1, 
/* out0446_had-eta6-phi22*/	5, 5, 0, 2, 5, 1, 12, 11, 0, 3, 12, 2, 9, 152, 0, 4, 
/* out0447_had-eta7-phi22*/	6, 4, 1, 3, 5, 1, 2, 5, 2, 1, 11, 0, 7, 11, 2, 9, 151, 0, 3, 
/* out0448_had-eta8-phi22*/	4, 4, 1, 5, 10, 0, 11, 11, 2, 3, 151, 0, 3, 
/* out0449_had-eta9-phi22*/	4, 3, 1, 1, 10, 0, 2, 10, 2, 12, 151, 0, 2, 
/* out0450_had-eta10-phi22*/	3, 9, 0, 11, 10, 2, 1, 150, 0, 6, 
/* out0451_had-eta11-phi22*/	4, 9, 0, 1, 9, 1, 2, 9, 2, 8, 150, 0, 2, 
/* out0452_had-eta12-phi22*/	2, 8, 0, 6, 9, 2, 3, 
/* out0453_had-eta13-phi22*/	3, 8, 0, 3, 8, 1, 3, 8, 2, 1, 
/* out0454_had-eta14-phi22*/	2, 8, 1, 2, 8, 2, 4, 
/* out0455_had-eta15-phi22*/	3, 7, 0, 3, 7, 1, 1, 8, 2, 1, 
/* out0456_had-eta16-phi22*/	2, 7, 0, 1, 7, 1, 4, 
/* out0457_had-eta17-phi22*/	1, 7, 1, 3, 
/* out0458_had-eta18-phi22*/	2, 7, 1, 1, 7, 2, 1, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	0, 
/* out0462_had-eta2-phi23*/	1, 154, 0, 6, 
/* out0463_had-eta3-phi23*/	2, 153, 0, 3, 154, 0, 2, 
/* out0464_had-eta4-phi23*/	3, 13, 0, 9, 13, 1, 3, 153, 0, 4, 
/* out0465_had-eta5-phi23*/	6, 12, 0, 8, 12, 1, 7, 13, 0, 7, 13, 1, 6, 152, 0, 4, 153, 0, 1, 
/* out0466_had-eta6-phi23*/	5, 11, 0, 3, 11, 1, 1, 12, 1, 9, 12, 2, 7, 152, 0, 4, 
/* out0467_had-eta7-phi23*/	4, 11, 0, 3, 11, 1, 14, 11, 2, 2, 151, 0, 3, 
/* out0468_had-eta8-phi23*/	5, 10, 0, 3, 10, 1, 5, 11, 1, 1, 11, 2, 2, 151, 0, 3, 
/* out0469_had-eta9-phi23*/	3, 10, 1, 11, 10, 2, 1, 151, 0, 2, 
/* out0470_had-eta10-phi23*/	4, 9, 0, 1, 9, 1, 5, 10, 2, 1, 150, 0, 6, 
/* out0471_had-eta11-phi23*/	2, 9, 1, 8, 150, 0, 2, 
/* out0472_had-eta12-phi23*/	3, 8, 1, 2, 9, 1, 1, 9, 2, 1, 
/* out0473_had-eta13-phi23*/	1, 8, 1, 6, 
/* out0474_had-eta14-phi23*/	1, 8, 1, 3, 
/* out0475_had-eta15-phi23*/	1, 7, 1, 1, 
/* out0476_had-eta16-phi23*/	1, 7, 1, 3, 
/* out0477_had-eta17-phi23*/	1, 7, 1, 3, 
/* out0478_had-eta18-phi23*/	0, 
/* out0479_had-eta19-phi23*/	0, 
};