parameter integer matrixH [0:8564] = {
/* num inputs = 190(in0-in189) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 12 */
//* total number of input in adders 2694 */

/* out0000_em-eta0-phi0*/	1,145,0,7,
/* out0001_em-eta1-phi0*/	2,145,0,9,145,1,9,
/* out0002_em-eta2-phi0*/	3,141,0,1,144,0,11,145,1,7,
/* out0003_em-eta3-phi0*/	7,140,0,15,140,1,1,141,0,10,141,1,12,141,2,16,144,0,5,144,1,12,
/* out0004_em-eta4-phi0*/	8,138,0,2,138,1,8,140,0,1,140,1,15,140,2,13,141,1,3,143,0,13,144,1,4,
/* out0005_em-eta5-phi0*/	6,137,0,5,137,1,16,137,2,6,140,2,3,143,0,3,143,1,14,
/* out0006_em-eta6-phi0*/	7,96,0,2,136,0,7,136,1,16,136,2,13,137,0,7,142,0,16,143,1,2,
/* out0007_em-eta7-phi0*/	6,95,1,6,95,2,1,96,0,1,136,0,9,136,2,3,142,1,16,
/* out0008_em-eta8-phi0*/	4,94,1,14,95,0,5,95,1,10,142,2,15,
/* out0009_em-eta9-phi0*/	7,94,1,1,94,2,10,95,0,3,47,0,13,47,1,12,47,2,2,142,2,1,
/* out0010_em-eta10-phi0*/	8,34,4,1,94,0,7,94,1,1,94,2,4,46,0,1,46,1,4,47,0,3,47,2,9,
/* out0011_em-eta11-phi0*/	9,34,1,9,34,2,2,34,4,2,35,0,2,35,1,15,94,0,2,46,0,6,46,1,6,46,2,2,
/* out0012_em-eta12-phi0*/	9,32,5,15,34,0,14,34,1,7,34,2,5,34,3,3,45,0,6,45,1,2,46,0,9,46,2,7,
/* out0013_em-eta13-phi0*/	9,32,5,1,33,0,15,33,2,3,33,4,2,33,5,15,34,0,2,34,3,2,45,0,5,45,1,5,
/* out0014_em-eta14-phi0*/	8,32,2,3,33,0,1,33,2,1,33,3,2,33,4,14,33,5,1,45,0,4,45,2,5,
/* out0015_em-eta15-phi0*/	8,32,0,3,32,1,16,32,2,13,32,3,9,44,0,7,44,1,4,45,0,1,45,2,2,
/* out0016_em-eta16-phi0*/	4,32,0,13,42,4,9,44,0,5,44,1,1,
/* out0017_em-eta17-phi0*/	4,42,4,7,43,1,5,44,0,3,44,2,2,
/* out0018_em-eta18-phi0*/	4,42,1,1,43,1,9,44,0,1,44,2,1,
/* out0019_em-eta19-phi0*/	1,42,1,3,
/* out0020_em-eta0-phi1*/	1,145,3,7,
/* out0021_em-eta1-phi1*/	2,145,2,9,145,3,9,
/* out0022_em-eta2-phi1*/	3,139,1,3,144,3,11,145,2,7,
/* out0023_em-eta3-phi1*/	9,138,1,1,138,2,2,139,0,16,139,1,10,139,2,4,141,0,5,141,1,1,144,2,12,144,3,5,
/* out0024_em-eta4-phi1*/	7,97,1,1,98,0,1,138,0,12,138,1,7,138,2,14,143,3,13,144,2,4,
/* out0025_em-eta5-phi1*/	7,97,0,10,97,1,5,137,0,2,137,2,10,138,0,2,143,2,14,143,3,3,
/* out0026_em-eta6-phi1*/	7,96,0,4,96,1,14,96,2,2,97,0,1,137,0,2,142,5,16,143,2,2,
/* out0027_em-eta7-phi1*/	6,95,2,6,96,0,9,96,2,4,107,0,1,107,1,1,142,4,16,
/* out0028_em-eta8-phi1*/	6,95,0,6,95,2,9,106,1,1,107,0,1,43,2,2,142,3,15,
/* out0029_em-eta9-phi1*/	10,94,2,1,95,0,2,106,1,10,42,0,1,42,1,2,43,1,4,43,2,11,47,1,4,47,2,2,142,3,1,
/* out0030_em-eta10-phi1*/	9,34,4,7,94,0,7,94,2,1,106,0,4,106,1,4,42,0,11,42,1,1,46,1,1,47,2,3,
/* out0031_em-eta11-phi1*/	11,34,4,6,34,5,11,35,0,14,35,1,1,35,4,4,35,5,1,41,0,1,42,0,3,42,2,1,46,1,5,46,2,3,
/* out0032_em-eta12-phi1*/	7,34,2,9,34,3,4,35,3,7,35,4,12,41,0,6,45,1,2,46,2,4,
/* out0033_em-eta13-phi1*/	8,33,2,7,34,3,7,35,3,6,44,1,3,45,1,3,41,0,2,45,1,7,45,2,1,
/* out0034_em-eta14-phi1*/	6,33,2,5,33,3,9,44,0,3,44,1,5,40,0,1,45,2,7,
/* out0035_em-eta15-phi1*/	8,32,3,7,33,3,5,42,5,4,43,5,1,44,0,2,40,0,1,44,1,5,45,2,1,
/* out0036_em-eta16-phi1*/	4,42,5,12,43,0,2,44,1,4,44,2,2,
/* out0037_em-eta17-phi1*/	3,43,0,11,43,1,1,44,2,5,
/* out0038_em-eta18-phi1*/	5,42,1,4,42,2,4,43,0,2,43,1,1,44,2,2,
/* out0039_em-eta19-phi1*/	2,42,0,2,42,1,6,
/* out0040_em-eta0-phi2*/	1,149,0,7,
/* out0041_em-eta1-phi2*/	2,149,0,9,149,1,9,
/* out0042_em-eta2-phi2*/	4,99,2,2,139,1,1,148,0,11,149,1,7,
/* out0043_em-eta3-phi2*/	8,98,1,10,99,0,8,99,1,16,99,2,4,139,1,2,139,2,12,148,0,5,148,1,12,
/* out0044_em-eta4-phi2*/	7,97,1,4,98,0,15,98,1,5,98,2,9,109,1,1,147,0,13,148,1,4,
/* out0045_em-eta5-phi2*/	7,97,0,3,97,1,6,97,2,15,108,1,1,109,1,2,147,0,3,147,1,14,
/* out0046_em-eta6-phi2*/	8,96,1,2,96,2,6,97,0,2,97,2,1,108,0,1,108,1,12,146,0,16,147,1,2,
/* out0047_em-eta7-phi2*/	5,96,2,4,107,0,1,107,1,12,108,0,2,146,1,16,
/* out0048_em-eta8-phi2*/	8,106,2,1,107,0,13,107,2,2,37,0,1,37,2,1,43,1,2,43,2,3,146,2,15,
/* out0049_em-eta9-phi2*/	6,106,1,1,106,2,11,37,2,9,42,1,5,43,1,10,146,2,1,
/* out0050_em-eta10-phi2*/	6,46,4,2,106,0,10,106,2,1,42,0,1,42,1,8,42,2,8,
/* out0051_em-eta11-phi2*/	8,34,5,5,35,2,1,35,5,13,46,4,12,47,1,4,106,0,1,41,1,7,42,2,6,
/* out0052_em-eta12-phi2*/	9,35,2,15,35,3,2,35,5,2,44,4,5,46,1,1,47,1,5,41,0,5,41,1,4,41,2,3,
/* out0053_em-eta13-phi2*/	8,35,3,1,44,1,1,44,4,5,45,0,5,45,1,13,40,1,2,41,0,2,41,2,4,
/* out0054_em-eta14-phi2*/	7,44,0,3,44,1,7,44,2,10,44,3,1,45,0,1,40,0,6,40,1,2,
/* out0055_em-eta15-phi2*/	4,43,5,5,44,0,8,44,3,5,40,0,6,
/* out0056_em-eta16-phi2*/	7,43,2,1,43,4,4,43,5,10,39,1,1,40,0,1,44,1,2,44,2,2,
/* out0057_em-eta17-phi2*/	5,42,2,3,43,0,1,43,4,9,39,1,2,44,2,2,
/* out0058_em-eta18-phi2*/	6,42,0,1,42,1,1,42,2,8,42,3,2,39,0,1,39,1,1,
/* out0059_em-eta19-phi2*/	2,42,0,9,42,1,1,
/* out0060_em-eta0-phi3*/	1,149,3,7,
/* out0061_em-eta1-phi3*/	2,149,2,9,149,3,9,
/* out0062_em-eta2-phi3*/	5,99,2,4,111,1,3,111,2,3,148,3,11,149,2,7,
/* out0063_em-eta3-phi3*/	9,98,1,1,98,2,1,99,0,8,99,2,6,110,1,11,110,2,7,111,2,10,148,2,12,148,3,5,
/* out0064_em-eta4-phi3*/	7,98,2,6,109,1,6,109,2,9,110,0,9,110,1,5,147,3,13,148,2,4,
/* out0065_em-eta5-phi3*/	7,108,2,4,109,0,14,109,1,7,109,2,3,119,1,1,147,2,14,147,3,3,
/* out0066_em-eta6-phi3*/	6,108,0,8,108,1,3,108,2,12,119,1,1,146,5,16,147,2,2,
/* out0067_em-eta7-phi3*/	5,107,1,3,107,2,4,108,0,5,118,1,7,146,4,16,
/* out0068_em-eta8-phi3*/	5,107,2,10,117,1,5,118,1,1,37,0,5,146,3,15,
/* out0069_em-eta9-phi3*/	7,106,2,2,117,0,8,117,1,3,37,0,9,37,1,9,37,2,5,146,3,1,
/* out0070_em-eta10-phi3*/	12,46,5,13,47,0,1,47,4,2,47,5,12,106,0,1,106,2,1,117,0,2,36,0,5,36,1,6,37,1,2,37,2,1,42,2,1,
/* out0071_em-eta11-phi3*/	9,46,2,7,46,4,2,46,5,3,47,0,15,47,1,5,47,4,5,36,0,11,36,2,1,41,1,2,
/* out0072_em-eta12-phi3*/	9,44,4,4,44,5,3,46,0,4,46,1,15,46,2,2,47,1,2,35,0,2,41,1,3,41,2,6,
/* out0073_em-eta13-phi3*/	8,44,4,2,44,5,11,45,0,9,45,4,3,45,5,2,35,0,3,40,1,4,41,2,3,
/* out0074_em-eta14-phi3*/	7,44,2,6,45,0,1,45,3,2,45,4,12,40,0,1,40,1,6,40,2,2,
/* out0075_em-eta15-phi3*/	4,43,2,1,44,3,10,45,3,6,40,2,6,
/* out0076_em-eta16-phi3*/	4,43,2,13,43,3,1,39,1,4,40,2,2,
/* out0077_em-eta17-phi3*/	3,43,3,9,43,4,3,39,1,4,
/* out0078_em-eta18-phi3*/	3,42,2,1,42,3,9,39,0,5,
/* out0079_em-eta19-phi3*/	3,0,0,3,42,0,4,42,3,2,
/* out0080_em-eta0-phi4*/	1,153,0,7,
/* out0081_em-eta1-phi4*/	2,153,0,9,153,1,9,
/* out0082_em-eta2-phi4*/	4,111,1,4,121,1,1,152,0,11,153,1,7,
/* out0083_em-eta3-phi4*/	7,110,2,9,111,1,9,111,2,3,121,0,12,121,1,12,152,0,5,152,1,12,
/* out0084_em-eta4-phi4*/	8,109,2,2,110,0,7,120,0,3,120,1,15,120,2,7,121,0,1,151,0,13,152,1,4,
/* out0085_em-eta5-phi4*/	8,109,0,2,109,2,2,119,1,8,119,2,9,120,0,5,120,1,1,151,0,3,151,1,14,
/* out0086_em-eta6-phi4*/	6,118,1,1,118,2,5,119,0,11,119,1,6,150,0,16,151,1,2,
/* out0087_em-eta7-phi4*/	4,118,0,6,118,1,7,118,2,7,150,1,16,
/* out0088_em-eta8-phi4*/	4,117,1,6,117,2,2,118,0,7,150,2,15,
/* out0089_em-eta9-phi4*/	8,117,0,3,117,1,2,117,2,9,37,0,1,37,1,5,38,0,7,38,2,11,150,2,1,
/* out0090_em-eta10-phi4*/	8,47,2,15,47,5,4,48,0,1,117,0,3,117,2,2,36,1,10,36,2,3,38,2,5,
/* out0091_em-eta11-phi4*/	7,46,2,6,46,3,8,47,2,1,47,3,14,47,4,9,35,1,1,36,2,12,
/* out0092_em-eta12-phi4*/	8,6,5,1,7,5,7,44,5,1,46,0,12,46,2,1,46,3,6,35,0,3,35,1,8,
/* out0093_em-eta13-phi4*/	7,6,4,2,6,5,8,44,5,1,45,2,1,45,5,12,35,0,7,35,2,2,
/* out0094_em-eta14-phi4*/	10,3,2,1,45,2,14,45,3,3,45,4,1,45,5,2,29,1,2,35,0,1,35,2,1,40,1,2,40,2,3,
/* out0095_em-eta15-phi4*/	6,3,2,2,3,5,10,45,2,1,45,3,5,29,1,3,40,2,3,
/* out0096_em-eta16-phi4*/	5,2,5,12,3,5,2,43,2,1,39,1,2,39,2,3,
/* out0097_em-eta17-phi4*/	6,2,4,6,2,5,1,43,3,5,39,0,2,39,1,2,39,2,3,
/* out0098_em-eta18-phi4*/	6,0,1,7,1,1,1,2,4,1,42,3,3,43,3,1,39,0,6,
/* out0099_em-eta19-phi4*/	2,0,0,9,0,1,3,
/* out0100_em-eta0-phi5*/	1,153,3,7,
/* out0101_em-eta1-phi5*/	2,153,2,9,153,3,9,
/* out0102_em-eta2-phi5*/	2,152,3,11,153,2,7,
/* out0103_em-eta3-phi5*/	5,121,0,2,121,1,3,121,2,16,152,2,12,152,3,5,
/* out0104_em-eta4-phi5*/	7,51,0,1,51,1,3,120,0,5,120,2,9,121,0,1,151,3,13,152,2,4,
/* out0105_em-eta5-phi5*/	7,51,0,15,51,1,1,51,2,3,119,2,6,120,0,3,151,2,14,151,3,3,
/* out0106_em-eta6-phi5*/	7,50,0,11,50,1,4,51,2,1,119,0,5,119,2,1,150,5,16,151,2,2,
/* out0107_em-eta7-phi5*/	7,49,0,1,49,1,3,50,0,5,50,2,4,118,0,2,118,2,4,150,4,16,
/* out0108_em-eta8-phi5*/	5,49,0,13,49,1,1,49,2,1,118,0,1,150,3,15,
/* out0109_em-eta9-phi5*/	8,48,0,2,48,1,3,49,0,2,49,2,3,117,2,3,38,0,9,38,1,10,150,3,1,
/* out0110_em-eta10-phi5*/	6,48,0,10,48,1,1,48,2,1,31,0,2,31,1,7,38,1,6,
/* out0111_em-eta11-phi5*/	7,7,2,8,46,3,2,47,3,2,48,0,3,48,2,3,31,0,13,35,1,1,
/* out0112_em-eta12-phi5*/	7,7,2,8,7,3,3,7,4,11,7,5,9,31,0,1,35,1,6,35,2,4,
/* out0113_em-eta13-phi5*/	6,6,4,4,6,5,7,7,0,12,7,1,2,29,2,1,35,2,9,
/* out0114_em-eta14-phi5*/	6,3,2,9,3,3,1,6,4,10,7,1,2,29,1,1,29,2,6,
/* out0115_em-eta15-phi5*/	5,3,2,4,3,3,3,3,4,8,3,5,4,29,1,7,
/* out0116_em-eta16-phi5*/	5,2,5,2,3,0,10,3,4,4,29,1,3,39,2,2,
/* out0117_em-eta17-phi5*/	5,2,4,6,2,5,1,3,0,2,3,1,3,39,2,5,
/* out0118_em-eta18-phi5*/	7,0,1,2,0,2,1,1,0,1,1,1,11,2,4,3,39,0,2,39,2,3,
/* out0119_em-eta19-phi5*/	5,0,0,4,0,1,4,0,2,11,0,3,2,1,0,3,
/* out0120_em-eta0-phi6*/	1,157,0,7,
/* out0121_em-eta1-phi6*/	2,157,0,9,157,1,9,
/* out0122_em-eta2-phi6*/	2,156,0,11,157,1,7,
/* out0123_em-eta3-phi6*/	5,60,0,16,60,1,3,60,2,2,156,0,5,156,1,12,
/* out0124_em-eta4-phi6*/	6,51,1,4,59,0,5,59,1,9,60,2,1,155,0,13,156,1,4,
/* out0125_em-eta5-phi6*/	7,51,1,8,51,2,11,58,0,5,58,1,1,59,0,3,155,0,3,155,1,14,
/* out0126_em-eta6-phi6*/	6,50,1,12,50,2,3,51,2,1,58,0,6,154,0,16,155,1,2,
/* out0127_em-eta7-phi6*/	5,49,1,4,50,2,9,57,0,2,57,1,4,154,1,16,
/* out0128_em-eta8-phi6*/	4,49,1,8,49,2,7,57,0,1,154,2,15,
/* out0129_em-eta9-phi6*/	7,48,1,5,49,2,5,56,0,3,33,0,11,33,1,2,33,2,10,154,2,1,
/* out0130_em-eta10-phi6*/	6,48,1,6,48,2,5,31,1,8,31,2,2,33,1,1,33,2,6,
/* out0131_em-eta11-phi6*/	8,6,3,2,7,3,7,18,5,2,19,5,2,48,2,6,30,2,1,31,1,1,31,2,13,
/* out0132_em-eta12-phi6*/	8,6,0,1,6,2,8,6,3,12,7,3,6,7,4,5,30,1,4,30,2,6,31,2,1,
/* out0133_em-eta13-phi6*/	6,6,1,9,6,2,8,7,0,4,7,1,3,29,2,1,30,1,9,
/* out0134_em-eta14-phi6*/	6,2,3,2,3,3,8,6,1,2,7,1,9,29,0,1,29,2,7,
/* out0135_em-eta15-phi6*/	5,2,2,5,2,3,5,3,3,4,3,4,4,29,0,6,
/* out0136_em-eta16-phi6*/	5,2,1,1,2,2,11,3,0,3,24,1,2,29,0,4,
/* out0137_em-eta17-phi6*/	4,2,1,2,3,0,1,3,1,9,24,1,4,
/* out0138_em-eta18-phi6*/	5,0,4,7,1,1,4,3,1,3,24,0,2,24,1,2,
/* out0139_em-eta19-phi6*/	6,0,2,4,0,3,6,0,5,1,1,0,11,1,3,1,1,5,1,
/* out0140_em-eta0-phi7*/	1,157,3,7,
/* out0141_em-eta1-phi7*/	2,157,2,9,157,3,9,
/* out0142_em-eta2-phi7*/	5,60,1,1,71,0,1,71,2,3,156,3,11,157,2,7,
/* out0143_em-eta3-phi7*/	6,60,1,12,60,2,12,70,1,9,71,0,11,156,2,12,156,3,5,
/* out0144_em-eta4-phi7*/	8,59,0,3,59,1,7,59,2,15,60,2,1,69,0,2,70,0,7,155,3,13,156,2,4,
/* out0145_em-eta5-phi7*/	8,58,0,2,58,1,15,58,2,1,59,0,5,59,2,1,69,0,4,155,2,14,155,3,3,
/* out0146_em-eta6-phi7*/	6,57,1,5,57,2,1,58,0,3,58,2,14,154,5,16,155,2,2,
/* out0147_em-eta7-phi7*/	4,57,0,6,57,1,7,57,2,7,154,4,16,
/* out0148_em-eta8-phi7*/	4,56,0,2,56,1,6,57,0,7,154,3,15,
/* out0149_em-eta9-phi7*/	8,56,0,9,56,1,2,56,2,3,33,0,5,33,1,10,34,0,2,34,2,5,154,3,1,
/* out0150_em-eta10-phi7*/	9,19,2,15,19,3,4,48,1,1,48,2,1,56,0,2,56,2,3,32,1,3,32,2,10,33,1,3,
/* out0151_em-eta11-phi7*/	7,18,5,8,19,0,6,19,2,1,19,4,9,19,5,14,30,2,1,32,1,12,
/* out0152_em-eta12-phi7*/	8,6,0,8,6,3,2,17,2,1,18,4,12,18,5,6,19,0,1,30,0,3,30,2,8,
/* out0153_em-eta13-phi7*/	6,6,0,7,6,1,4,17,2,9,17,5,7,30,0,7,30,1,2,
/* out0154_em-eta14-phi7*/	10,2,3,2,6,1,1,16,5,10,17,5,8,25,1,3,25,2,2,29,0,2,29,2,1,30,0,1,30,1,1,
/* out0155_em-eta15-phi7*/	6,2,0,6,2,3,7,16,4,3,16,5,3,25,1,3,29,0,3,
/* out0156_em-eta16-phi7*/	5,2,0,9,2,1,5,5,2,1,24,1,4,24,2,2,
/* out0157_em-eta17-phi7*/	4,2,1,8,5,5,5,24,0,1,24,1,4,
/* out0158_em-eta18-phi7*/	5,0,4,8,3,1,1,4,5,3,5,5,1,24,0,5,
/* out0159_em-eta19-phi7*/	6,0,3,4,0,4,1,0,5,11,1,0,1,1,3,7,1,5,7,
/* out0160_em-eta0-phi8*/	1,161,0,7,
/* out0161_em-eta1-phi8*/	2,161,0,9,161,1,9,
/* out0162_em-eta2-phi8*/	5,71,2,7,82,0,4,82,1,2,160,0,11,161,1,7,
/* out0163_em-eta3-phi8*/	11,70,1,7,70,2,11,71,0,4,71,2,6,81,0,1,81,1,1,82,0,12,82,1,1,82,2,9,160,0,5,160,1,12,
/* out0164_em-eta4-phi8*/	7,69,0,2,69,1,13,70,0,9,70,2,5,81,0,6,159,0,13,160,1,4,
/* out0165_em-eta5-phi8*/	6,68,1,4,69,0,8,69,1,2,69,2,14,159,0,3,159,1,14,
/* out0166_em-eta6-phi8*/	6,58,2,1,68,0,8,68,1,12,68,2,3,158,0,16,159,1,2,
/* out0167_em-eta7-phi8*/	4,57,2,7,67,1,8,68,0,5,158,1,16,
/* out0168_em-eta8-phi8*/	6,56,1,5,57,2,1,67,0,7,67,1,3,34,0,4,158,2,15,
/* out0169_em-eta9-phi8*/	7,56,1,3,56,2,8,66,1,2,34,0,9,34,1,7,34,2,8,158,2,1,
/* out0170_em-eta10-phi8*/	12,18,2,1,18,3,13,19,3,12,19,4,2,56,2,2,66,0,1,66,1,1,27,1,1,32,0,5,32,2,6,34,1,1,34,2,3,
/* out0171_em-eta11-phi8*/	9,18,0,2,18,1,5,18,2,15,18,3,3,19,0,7,19,4,5,26,2,2,32,0,11,32,1,1,
/* out0172_em-eta12-phi8*/	9,17,2,2,17,3,5,18,1,2,18,4,4,19,0,2,19,1,15,26,1,6,26,2,3,30,0,2,
/* out0173_em-eta13-phi8*/	8,16,2,1,17,2,4,17,3,9,17,4,11,17,5,1,25,2,4,26,1,3,30,0,3,
/* out0174_em-eta14-phi8*/	7,16,2,1,16,5,2,17,0,13,17,4,5,25,0,1,25,1,2,25,2,6,
/* out0175_em-eta15-phi8*/	5,5,2,1,16,4,13,16,5,1,17,1,3,25,1,6,
/* out0176_em-eta16-phi8*/	5,2,0,1,5,2,13,5,5,1,24,2,5,25,1,2,
/* out0177_em-eta17-phi8*/	4,5,4,3,5,5,9,24,0,2,24,2,4,
/* out0178_em-eta18-phi8*/	3,4,5,9,5,0,1,24,0,5,
/* out0179_em-eta19-phi8*/	6,0,3,4,0,5,4,1,3,8,1,5,8,4,4,4,4,5,2,
/* out0180_em-eta0-phi9*/	1,161,3,7,
/* out0181_em-eta1-phi9*/	2,161,2,9,161,3,9,
/* out0182_em-eta2-phi9*/	4,82,1,2,124,1,1,160,3,11,161,2,7,
/* out0183_em-eta3-phi9*/	7,81,1,10,82,1,11,82,2,7,124,0,5,124,1,9,160,2,12,160,3,5,
/* out0184_em-eta4-phi9*/	7,69,1,1,80,1,4,81,0,9,81,1,5,81,2,15,159,3,13,160,2,4,
/* out0185_em-eta5-phi9*/	7,68,2,1,69,2,2,80,0,15,80,1,6,80,2,3,159,2,14,159,3,3,
/* out0186_em-eta6-phi9*/	7,68,0,1,68,2,12,79,1,8,80,0,1,80,2,2,158,5,16,159,2,2,
/* out0187_em-eta7-phi9*/	5,67,1,5,67,2,8,68,0,2,79,0,4,158,4,16,
/* out0188_em-eta8-phi9*/	8,66,1,1,67,0,9,67,2,6,28,0,3,28,1,2,34,0,1,34,1,1,158,3,15,
/* out0189_em-eta9-phi9*/	6,66,1,11,66,2,1,27,2,5,28,1,10,34,1,7,158,3,1,
/* out0190_em-eta10-phi9*/	6,18,0,2,66,0,10,66,1,1,27,0,1,27,1,8,27,2,8,
/* out0191_em-eta11-phi9*/	8,18,0,12,18,1,4,20,3,5,21,2,1,21,3,13,66,0,1,26,2,7,27,1,6,
/* out0192_em-eta12-phi9*/	10,16,3,3,17,3,2,18,1,5,19,1,1,21,2,15,21,3,2,21,5,2,26,0,5,26,1,3,26,2,4,
/* out0193_em-eta13-phi9*/	7,16,0,6,16,2,6,16,3,13,21,5,1,25,2,2,26,0,2,26,1,4,
/* out0194_em-eta14-phi9*/	7,16,0,1,16,1,9,16,2,8,17,0,3,17,1,1,25,0,6,25,2,2,
/* out0195_em-eta15-phi9*/	4,5,3,5,16,1,1,17,1,12,25,0,6,
/* out0196_em-eta16-phi9*/	7,5,2,1,5,3,10,5,4,4,20,1,2,20,2,2,24,2,1,25,0,1,
/* out0197_em-eta17-phi9*/	5,4,2,1,5,0,3,5,4,9,20,1,2,24,2,3,
/* out0198_em-eta18-phi9*/	6,4,4,1,4,5,2,5,0,8,5,1,1,24,0,1,24,2,1,
/* out0199_em-eta19-phi9*/	2,4,4,9,5,1,1,
/* out0200_em-eta0-phi10*/	1,165,0,7,
/* out0201_em-eta1-phi10*/	2,165,0,9,165,1,9,
/* out0202_em-eta2-phi10*/	4,124,1,2,124,2,2,164,0,11,165,1,7,
/* out0203_em-eta3-phi10*/	9,123,1,2,123,2,1,124,0,11,124,1,4,124,2,14,125,0,2,125,2,6,164,0,5,164,1,12,
/* out0204_em-eta4-phi10*/	7,80,1,1,81,2,1,123,0,12,123,1,14,123,2,7,163,0,13,164,1,4,
/* out0205_em-eta5-phi10*/	7,80,1,5,80,2,10,122,0,9,122,1,3,123,0,2,163,0,3,163,1,14,
/* out0206_em-eta6-phi10*/	7,79,0,1,79,1,8,79,2,11,80,2,1,122,0,2,162,0,16,163,1,2,
/* out0207_em-eta7-phi10*/	5,67,2,1,78,1,6,79,0,11,79,2,2,162,1,16,
/* out0208_em-eta8-phi10*/	6,66,2,1,67,2,1,78,0,6,78,1,9,28,0,2,162,2,15,
/* out0209_em-eta9-phi10*/	9,66,2,10,78,0,2,23,1,2,23,2,4,27,0,1,27,2,2,28,0,11,28,1,4,162,2,1,
/* out0210_em-eta10-phi10*/	8,20,0,6,66,0,4,66,2,4,88,1,1,22,2,1,23,1,3,27,0,11,27,2,1,
/* out0211_em-eta11-phi10*/	11,20,0,7,20,1,1,20,2,14,20,3,11,21,3,1,21,4,4,22,1,3,22,2,5,26,0,1,27,0,3,27,1,1,
/* out0212_em-eta12-phi10*/	7,20,5,3,21,0,8,21,4,12,21,5,6,21,2,2,22,1,4,26,0,6,
/* out0213_em-eta13-phi10*/	8,16,0,6,20,5,7,21,5,7,28,5,2,29,5,3,21,1,1,21,2,7,26,0,2,
/* out0214_em-eta14-phi10*/	6,16,0,3,16,1,4,28,4,3,28,5,9,21,1,7,25,0,1,
/* out0215_em-eta15-phi10*/	7,4,3,4,5,3,1,16,1,2,28,4,10,20,2,5,21,1,1,25,0,1,
/* out0216_em-eta16-phi10*/	4,4,2,2,4,3,12,20,1,2,20,2,4,
/* out0217_em-eta17-phi10*/	3,4,1,1,4,2,11,20,1,5,
/* out0218_em-eta18-phi10*/	5,4,1,1,4,2,2,5,0,4,5,1,4,20,1,2,
/* out0219_em-eta19-phi10*/	2,4,4,2,5,1,6,
/* out0220_em-eta0-phi11*/	1,165,3,7,
/* out0221_em-eta1-phi11*/	2,165,2,9,165,3,9,
/* out0222_em-eta2-phi11*/	3,125,0,1,164,3,11,165,2,7,
/* out0223_em-eta3-phi11*/	6,125,0,13,125,1,15,125,2,9,132,1,1,164,2,12,164,3,5,
/* out0224_em-eta4-phi11*/	9,122,1,1,123,0,2,123,2,8,125,1,1,125,2,1,132,0,14,132,1,7,163,3,13,164,2,4,
/* out0225_em-eta5-phi11*/	6,122,0,3,122,1,12,122,2,11,132,0,2,163,2,14,163,3,3,
/* out0226_em-eta6-phi11*/	6,79,2,2,122,0,2,122,2,5,130,2,13,162,5,16,163,2,2,
/* out0227_em-eta7-phi11*/	6,78,1,1,78,2,6,79,2,1,130,1,8,130,2,3,162,4,16,
/* out0228_em-eta8-phi11*/	3,78,0,5,78,2,10,162,3,15,
/* out0229_em-eta9-phi11*/	7,78,0,3,88,1,3,88,2,8,23,0,5,23,1,2,23,2,12,162,3,1,
/* out0230_em-eta10-phi11*/	5,20,0,1,88,1,11,22,2,4,23,0,3,23,1,9,
/* out0231_em-eta11-phi11*/	9,20,0,2,20,1,15,20,2,2,21,0,2,21,1,9,88,1,1,22,0,6,22,1,2,22,2,6,
/* out0232_em-eta12-phi11*/	7,20,4,14,20,5,4,21,0,6,21,1,7,21,2,2,22,0,2,22,1,7,
/* out0233_em-eta13-phi11*/	7,20,4,2,20,5,2,29,2,7,29,4,1,29,5,12,21,0,5,21,2,5,
/* out0234_em-eta14-phi11*/	6,28,5,5,29,0,10,29,4,6,29,5,1,21,0,4,21,1,5,
/* out0235_em-eta15-phi11*/	6,28,4,3,29,0,5,29,1,10,20,0,1,20,2,4,21,1,2,
/* out0236_em-eta16-phi11*/	4,4,0,9,29,1,5,20,0,4,20,2,1,
/* out0237_em-eta17-phi11*/	4,4,0,7,4,1,5,20,0,3,20,1,2,
/* out0238_em-eta18-phi11*/	3,4,1,9,5,1,1,20,1,1,
/* out0239_em-eta19-phi11*/	1,5,1,3,
/* out0240_em-eta0-phi12*/	1,169,0,7,
/* out0241_em-eta1-phi12*/	2,169,0,9,169,1,9,
/* out0242_em-eta2-phi12*/	2,168,0,11,169,1,7,
/* out0243_em-eta3-phi12*/	6,132,1,1,134,0,15,134,1,9,134,2,13,168,0,5,168,1,12,
/* out0244_em-eta4-phi12*/	9,131,2,1,132,1,7,132,2,14,133,1,8,133,2,2,134,1,1,134,2,3,167,0,13,168,1,4,
/* out0245_em-eta5-phi12*/	6,131,0,3,131,1,11,131,2,12,132,2,2,167,0,3,167,1,14,
/* out0246_em-eta6-phi12*/	6,90,1,2,130,0,13,131,0,2,131,1,5,166,0,16,167,1,2,
/* out0247_em-eta7-phi12*/	5,89,2,7,90,1,1,130,0,3,130,1,8,166,1,16,
/* out0248_em-eta8-phi12*/	3,89,1,13,89,2,3,166,2,15,
/* out0249_em-eta9-phi12*/	8,88,0,2,88,2,8,89,1,3,18,1,1,19,0,13,19,2,4,23,0,5,166,2,1,
/* out0250_em-eta10-phi12*/	5,31,3,1,88,0,10,18,0,12,18,1,2,23,0,3,
/* out0251_em-eta11-phi12*/	10,31,2,15,31,3,9,31,4,4,31,5,2,88,0,2,17,0,1,17,1,1,18,0,4,18,2,2,22,0,6,
/* out0252_em-eta12-phi12*/	7,30,5,9,31,0,1,31,2,1,31,4,4,31,5,14,17,0,9,22,0,2,
/* out0253_em-eta13-phi12*/	8,29,2,9,29,3,11,29,4,2,30,4,1,30,5,4,17,0,4,17,2,1,21,0,4,
/* out0254_em-eta14-phi12*/	6,28,2,10,28,3,3,29,3,1,29,4,7,16,0,4,21,0,3,
/* out0255_em-eta15-phi12*/	6,28,0,1,28,1,10,28,2,6,29,0,1,16,0,6,20,0,1,
/* out0256_em-eta16-phi12*/	6,28,1,6,29,1,1,36,5,1,37,5,7,16,0,1,20,0,4,
/* out0257_em-eta17-phi12*/	3,36,5,11,15,0,3,20,0,3,
/* out0258_em-eta18-phi12*/	4,36,4,9,36,5,2,15,0,2,15,1,1,
/* out0259_em-eta19-phi12*/	1,36,4,4,
/* out0260_em-eta0-phi13*/	1,169,3,7,
/* out0261_em-eta1-phi13*/	2,169,2,9,169,3,9,
/* out0262_em-eta2-phi13*/	3,135,2,3,168,3,11,169,2,7,
/* out0263_em-eta3-phi13*/	8,133,2,4,134,0,1,134,1,6,135,0,4,135,1,16,135,2,10,168,2,12,168,3,5,
/* out0264_em-eta4-phi13*/	7,91,2,1,92,1,1,133,0,15,133,1,7,133,2,10,167,3,13,168,2,4,
/* out0265_em-eta5-phi13*/	8,91,1,2,91,2,12,131,0,9,131,2,3,133,0,1,133,1,1,167,2,14,167,3,3,
/* out0266_em-eta6-phi13*/	7,90,0,2,90,1,4,90,2,14,91,1,1,131,0,2,166,5,16,167,2,2,
/* out0267_em-eta7-phi13*/	7,89,0,1,89,2,5,90,0,4,90,1,9,101,1,1,101,2,1,166,4,16,
/* out0268_em-eta8-phi13*/	6,89,0,13,89,2,1,100,2,1,101,1,1,19,0,1,166,3,15,
/* out0269_em-eta9-phi13*/	8,88,0,1,89,0,2,100,2,10,14,0,7,18,1,3,19,0,2,19,2,12,166,3,1,
/* out0270_em-eta10-phi13*/	8,30,3,4,31,3,2,88,0,1,100,1,4,100,2,4,14,0,1,18,1,10,18,2,5,
/* out0271_em-eta11-phi13*/	9,30,0,3,30,1,1,30,2,12,30,3,12,31,3,4,31,4,6,12,0,1,17,1,5,18,2,8,
/* out0272_em-eta12-phi13*/	9,30,2,4,30,4,2,30,5,3,31,0,15,31,1,5,31,4,2,17,0,2,17,1,7,17,2,3,
/* out0273_em-eta13-phi13*/	7,28,3,2,29,3,4,30,4,13,38,5,3,39,5,3,16,1,1,17,2,8,
/* out0274_em-eta14-phi13*/	6,28,0,4,28,3,11,38,4,3,38,5,5,16,0,1,16,1,7,
/* out0275_em-eta15-phi13*/	6,28,0,11,37,2,5,38,4,2,16,0,3,16,1,1,16,2,3,
/* out0276_em-eta16-phi13*/	6,37,2,5,37,4,2,37,5,8,15,0,2,16,0,1,16,2,3,
/* out0277_em-eta17-phi13*/	5,36,5,1,37,0,6,37,4,4,37,5,1,15,0,6,
/* out0278_em-eta18-phi13*/	5,36,4,1,36,5,1,37,0,6,37,1,3,15,1,2,
/* out0279_em-eta19-phi13*/	2,36,4,2,37,1,6,
/* out0280_em-eta0-phi14*/	1,173,0,7,
/* out0281_em-eta1-phi14*/	2,173,0,9,173,1,9,
/* out0282_em-eta2-phi14*/	4,93,0,4,135,2,1,172,0,11,173,1,7,
/* out0283_em-eta3-phi14*/	8,92,2,10,93,0,7,93,1,1,93,2,15,135,0,12,135,2,2,172,0,5,172,1,12,
/* out0284_em-eta4-phi14*/	8,91,0,3,91,2,1,92,0,9,92,1,15,92,2,5,103,2,1,171,0,13,172,1,4,
/* out0285_em-eta5-phi14*/	7,91,0,13,91,1,10,91,2,2,102,2,1,103,2,2,171,0,3,171,1,14,
/* out0286_em-eta6-phi14*/	7,90,0,6,90,2,2,91,1,3,102,1,1,102,2,12,170,0,16,171,1,2,
/* out0287_em-eta7-phi14*/	5,90,0,4,101,1,1,101,2,12,102,1,2,170,1,16,
/* out0288_em-eta8-phi14*/	5,100,0,1,101,0,2,101,1,13,14,1,5,170,2,15,
/* out0289_em-eta9-phi14*/	6,100,0,11,100,2,1,14,0,6,14,1,9,14,2,5,170,2,1,
/* out0290_em-eta10-phi14*/	8,41,2,2,100,0,1,100,1,10,12,0,2,12,1,6,14,0,2,14,2,6,18,2,1,
/* out0291_em-eta11-phi14*/	8,30,0,13,30,1,5,41,2,13,41,5,4,100,1,1,12,0,11,12,1,1,12,2,1,
/* out0292_em-eta12-phi14*/	11,30,1,10,31,1,10,39,2,5,40,5,1,41,5,5,10,0,2,10,1,1,12,0,2,12,2,2,17,1,3,17,2,2,
/* out0293_em-eta13-phi14*/	8,31,1,1,38,5,1,39,2,5,39,4,5,39,5,13,10,0,7,16,1,1,17,2,2,
/* out0294_em-eta14-phi14*/	7,38,4,3,38,5,7,39,0,10,39,1,1,39,4,1,10,0,1,16,1,6,
/* out0295_em-eta15-phi14*/	5,37,2,4,37,3,1,38,4,8,39,1,5,16,2,6,
/* out0296_em-eta16-phi14*/	7,37,2,2,37,3,8,37,4,5,9,0,1,15,0,2,15,1,1,16,2,3,
/* out0297_em-eta17-phi14*/	5,36,2,7,37,0,1,37,4,5,15,0,1,15,1,5,
/* out0298_em-eta18-phi14*/	5,36,1,2,36,2,5,37,0,3,37,1,1,15,1,1,
/* out0299_em-eta19-phi14*/	2,36,1,4,37,1,6,
/* out0300_em-eta0-phi15*/	1,173,3,7,
/* out0301_em-eta1-phi15*/	2,173,2,9,173,3,9,
/* out0302_em-eta2-phi15*/	6,93,0,4,93,1,2,105,0,3,105,1,3,172,3,11,173,2,7,
/* out0303_em-eta3-phi15*/	10,92,0,1,92,2,1,93,0,1,93,1,13,93,2,1,104,0,7,104,2,11,105,1,10,172,2,12,172,3,5,
/* out0304_em-eta4-phi15*/	7,92,0,6,103,0,9,103,2,6,104,1,9,104,2,5,171,3,13,172,2,4,
/* out0305_em-eta5-phi15*/	6,102,0,4,103,0,3,103,1,14,103,2,7,171,2,14,171,3,3,
/* out0306_em-eta6-phi15*/	6,102,0,12,102,1,8,102,2,3,114,1,1,170,5,16,171,2,2,
/* out0307_em-eta7-phi15*/	6,101,0,4,101,2,3,102,1,5,113,1,4,113,2,3,170,4,16,
/* out0308_em-eta8-phi15*/	4,101,0,10,112,2,5,113,1,1,170,3,15,
/* out0309_em-eta9-phi15*/	8,100,0,2,112,1,8,112,2,3,13,1,5,13,2,4,14,1,2,14,2,4,170,3,1,
/* out0310_em-eta10-phi15*/	10,40,2,2,40,3,12,41,3,13,41,4,1,100,0,1,100,1,1,112,1,2,12,1,6,13,1,9,14,2,1,
/* out0311_em-eta11-phi15*/	9,40,2,5,41,0,7,41,2,1,41,3,3,41,4,15,41,5,5,11,1,1,12,1,3,12,2,10,
/* out0312_em-eta12-phi15*/	8,39,2,4,39,3,3,40,4,4,40,5,15,41,0,2,41,5,2,10,1,8,12,2,3,
/* out0313_em-eta13-phi15*/	8,38,2,3,38,3,2,39,2,2,39,3,11,39,4,9,10,0,4,10,1,3,10,2,3,
/* out0314_em-eta14-phi15*/	7,38,1,2,38,2,12,39,0,6,39,4,1,9,1,2,10,0,2,10,2,4,
/* out0315_em-eta15-phi15*/	6,37,3,1,38,1,6,39,1,10,9,0,5,9,1,1,16,2,1,
/* out0316_em-eta16-phi15*/	4,36,3,8,37,3,6,9,0,5,15,1,1,
/* out0317_em-eta17-phi15*/	5,36,0,2,36,2,3,36,3,7,9,0,1,15,1,5,
/* out0318_em-eta18-phi15*/	3,36,0,5,36,1,5,36,2,1,
/* out0319_em-eta19-phi15*/	5,8,3,3,8,5,1,9,3,2,9,5,2,36,1,5,
/* out0320_em-eta0-phi16*/	1,177,0,7,
/* out0321_em-eta1-phi16*/	2,177,0,9,177,1,9,
/* out0322_em-eta2-phi16*/	4,105,0,4,116,2,1,176,0,11,177,1,7,
/* out0323_em-eta3-phi16*/	7,104,0,9,105,0,9,105,1,3,116,1,12,116,2,12,176,0,5,176,1,12,
/* out0324_em-eta4-phi16*/	8,103,0,2,104,1,7,115,0,7,115,1,3,115,2,15,116,1,1,175,0,13,176,1,4,
/* out0325_em-eta5-phi16*/	9,103,0,2,103,1,2,114,0,2,114,1,1,114,2,15,115,1,5,115,2,1,175,0,3,175,1,14,
/* out0326_em-eta6-phi16*/	5,113,2,6,114,0,3,114,1,14,174,0,16,175,1,2,
/* out0327_em-eta7-phi16*/	4,113,0,7,113,1,5,113,2,7,174,1,16,
/* out0328_em-eta8-phi16*/	5,112,0,2,112,2,6,113,0,2,113,1,6,174,2,15,
/* out0329_em-eta9-phi16*/	6,112,0,9,112,1,3,112,2,2,13,0,3,13,2,12,174,2,1,
/* out0330_em-eta10-phi16*/	8,40,0,15,40,3,4,52,0,1,112,0,2,112,1,3,11,2,3,13,0,12,13,1,2,
/* out0331_em-eta11-phi16*/	7,40,0,1,40,1,14,40,2,9,41,0,6,41,1,8,11,1,8,11,2,5,
/* out0332_em-eta12-phi16*/	9,14,5,1,15,5,7,39,3,1,40,4,12,41,0,1,41,1,6,10,1,3,11,0,2,11,1,7,
/* out0333_em-eta13-phi16*/	8,14,4,2,14,5,8,38,0,1,38,3,12,39,3,1,10,1,1,10,2,6,48,1,2,
/* out0334_em-eta14-phi16*/	8,13,3,1,38,0,14,38,1,3,38,2,1,38,3,2,9,1,4,10,2,3,48,1,1,
/* out0335_em-eta15-phi16*/	7,13,2,6,13,3,6,38,0,1,38,1,5,9,0,1,9,1,5,9,2,1,
/* out0336_em-eta16-phi16*/	4,13,2,10,13,5,4,9,0,2,9,2,3,
/* out0337_em-eta17-phi16*/	5,13,5,7,36,0,4,36,3,1,9,0,1,9,2,2,
/* out0338_em-eta18-phi16*/	3,8,0,7,12,5,1,36,0,5,
/* out0339_em-eta19-phi16*/	6,8,0,1,8,2,1,8,3,11,8,5,7,9,3,13,9,5,13,
/* out0340_em-eta0-phi17*/	1,177,3,7,
/* out0341_em-eta1-phi17*/	2,177,2,9,177,3,9,
/* out0342_em-eta2-phi17*/	2,176,3,11,177,2,7,
/* out0343_em-eta3-phi17*/	5,116,0,16,116,1,2,116,2,3,176,2,12,176,3,5,
/* out0344_em-eta4-phi17*/	7,55,0,1,55,1,3,115,0,9,115,1,5,116,1,1,175,3,13,176,2,4,
/* out0345_em-eta5-phi17*/	8,55,0,15,55,1,1,55,2,3,114,0,5,114,2,1,115,1,3,175,2,14,175,3,3,
/* out0346_em-eta6-phi17*/	6,54,0,11,54,1,4,55,2,1,114,0,6,174,5,16,175,2,2,
/* out0347_em-eta7-phi17*/	5,53,1,4,54,0,5,54,2,4,113,0,6,174,4,16,
/* out0348_em-eta8-phi17*/	4,53,0,7,53,1,8,113,0,1,174,3,15,
/* out0349_em-eta9-phi17*/	8,52,0,2,52,1,3,53,0,5,112,0,3,13,0,1,51,0,3,51,1,8,174,3,1,
/* out0350_em-eta10-phi17*/	5,52,0,10,52,1,1,52,2,1,11,2,2,51,0,13,
/* out0351_em-eta11-phi17*/	7,15,2,8,40,1,2,41,1,2,52,0,3,52,2,3,11,0,7,11,2,6,
/* out0352_em-eta12-phi17*/	6,15,2,8,15,3,3,15,4,11,15,5,9,11,0,7,48,2,4,
/* out0353_em-eta13-phi17*/	6,14,4,4,14,5,7,15,0,12,15,1,2,48,1,6,48,2,4,
/* out0354_em-eta14-phi17*/	6,12,3,8,13,3,2,14,4,10,15,1,2,9,1,1,48,1,7,
/* out0355_em-eta15-phi17*/	6,12,2,3,12,3,4,13,3,7,13,4,5,9,1,3,9,2,4,
/* out0356_em-eta16-phi17*/	4,13,0,2,13,4,11,13,5,2,9,2,5,
/* out0357_em-eta17-phi17*/	4,12,5,8,13,0,2,13,5,3,9,2,1,
/* out0358_em-eta18-phi17*/	3,8,0,8,8,1,3,12,5,3,
/* out0359_em-eta19-phi17*/	6,8,2,11,8,3,2,8,5,6,9,0,4,9,3,1,9,5,1,
/* out0360_em-eta0-phi18*/	1,181,0,7,
/* out0361_em-eta1-phi18*/	2,181,0,9,181,1,9,
/* out0362_em-eta2-phi18*/	2,180,0,11,181,1,7,
/* out0363_em-eta3-phi18*/	4,65,0,9,65,1,11,180,0,5,180,1,12,
/* out0364_em-eta4-phi18*/	6,55,1,4,64,0,12,64,1,2,65,0,1,179,0,13,180,1,4,
/* out0365_em-eta5-phi18*/	8,55,1,8,55,2,11,63,0,5,63,1,1,64,0,2,64,2,1,179,0,3,179,1,14,
/* out0366_em-eta6-phi18*/	6,54,1,12,54,2,3,55,2,1,63,0,6,178,0,16,179,1,2,
/* out0367_em-eta7-phi18*/	5,53,1,3,53,2,2,54,2,9,62,0,6,178,1,16,
/* out0368_em-eta8-phi18*/	5,53,0,1,53,1,1,53,2,12,62,0,1,178,2,15,
/* out0369_em-eta9-phi18*/	9,52,1,5,53,0,3,53,2,2,61,0,1,61,1,2,50,1,1,51,1,8,51,2,3,178,2,1,
/* out0370_em-eta10-phi18*/	4,52,1,6,52,2,5,49,2,2,51,2,13,
/* out0371_em-eta11-phi18*/	7,14,3,2,15,3,7,26,5,2,27,5,2,52,2,6,49,1,7,49,2,6,
/* out0372_em-eta12-phi18*/	7,14,0,1,14,2,8,14,3,12,15,3,6,15,4,5,48,2,4,49,1,7,
/* out0373_em-eta13-phi18*/	6,14,1,9,14,2,8,15,0,4,15,1,3,48,0,6,48,2,4,
/* out0374_em-eta14-phi18*/	6,12,0,8,12,3,1,14,1,2,15,1,9,5,2,1,48,0,7,
/* out0375_em-eta15-phi18*/	6,12,0,4,12,1,3,12,2,9,12,3,3,5,1,4,5,2,3,
/* out0376_em-eta16-phi18*/	4,12,2,4,13,0,10,13,1,1,5,1,5,
/* out0377_em-eta17-phi18*/	5,12,4,6,12,5,4,13,0,2,13,1,1,5,1,1,
/* out0378_em-eta18-phi18*/	4,8,1,12,8,2,1,9,1,2,12,4,3,
/* out0379_em-eta19-phi18*/	5,8,2,3,8,4,4,8,5,2,9,0,12,9,1,3,
/* out0380_em-eta0-phi19*/	1,181,3,7,
/* out0381_em-eta1-phi19*/	2,181,2,9,181,3,9,
/* out0382_em-eta2-phi19*/	4,65,1,1,77,0,4,180,3,11,181,2,7,
/* out0383_em-eta3-phi19*/	8,65,0,5,65,1,4,65,2,16,76,1,9,77,0,9,77,2,3,180,2,12,180,3,5,
/* out0384_em-eta4-phi19*/	8,64,0,2,64,1,14,64,2,9,65,0,1,75,0,2,76,0,7,179,3,13,180,2,4,
/* out0385_em-eta5-phi19*/	7,63,0,2,63,1,15,63,2,1,64,2,6,75,0,4,179,2,14,179,3,3,
/* out0386_em-eta6-phi19*/	6,62,1,6,63,0,3,63,2,14,74,0,1,178,5,16,179,2,2,
/* out0387_em-eta7-phi19*/	4,62,0,7,62,1,7,62,2,5,178,4,16,
/* out0388_em-eta8-phi19*/	4,61,1,8,62,0,2,62,2,6,178,3,15,
/* out0389_em-eta9-phi19*/	6,61,0,8,61,1,5,61,2,1,50,1,3,50,2,12,178,3,1,
/* out0390_em-eta10-phi19*/	8,27,2,15,27,3,4,52,1,1,52,2,1,61,0,4,49,2,3,50,0,2,50,1,12,
/* out0391_em-eta11-phi19*/	7,26,5,8,27,0,6,27,2,1,27,4,9,27,5,14,49,0,8,49,2,5,
/* out0392_em-eta12-phi19*/	9,14,0,8,14,3,2,23,2,1,26,4,12,26,5,6,27,0,1,6,2,3,49,0,7,49,1,2,
/* out0393_em-eta13-phi19*/	7,14,0,7,14,1,4,23,2,9,23,5,7,6,1,6,6,2,1,48,0,2,
/* out0394_em-eta14-phi19*/	7,12,0,2,14,1,1,22,5,10,23,5,8,5,2,4,6,1,3,48,0,1,
/* out0395_em-eta15-phi19*/	7,12,0,2,12,1,11,22,4,3,22,5,3,5,0,1,5,1,1,5,2,5,
/* out0396_em-eta16-phi19*/	4,12,1,2,13,1,12,5,0,2,5,1,3,
/* out0397_em-eta17-phi19*/	6,11,2,4,11,3,1,12,4,6,13,1,1,5,0,1,5,1,2,
/* out0398_em-eta18-phi19*/	4,8,1,1,9,1,8,11,2,5,12,4,1,
/* out0399_em-eta19-phi19*/	2,8,4,8,9,1,3,
/* out0400_em-eta0-phi20*/	1,185,0,7,
/* out0401_em-eta1-phi20*/	2,185,0,9,185,1,9,
/* out0402_em-eta2-phi20*/	6,77,0,3,77,2,3,87,0,5,87,2,2,184,0,11,185,1,7,
/* out0403_em-eta3-phi20*/	9,76,1,7,76,2,11,77,2,10,86,1,1,87,0,2,87,1,2,87,2,14,184,0,5,184,1,12,
/* out0404_em-eta4-phi20*/	8,75,0,2,75,1,13,76,0,9,76,2,5,86,0,2,86,1,4,183,0,13,184,1,4,
/* out0405_em-eta5-phi20*/	6,74,1,4,75,0,8,75,1,2,75,2,14,183,0,3,183,1,14,
/* out0406_em-eta6-phi20*/	6,63,2,1,74,0,13,74,1,6,74,2,3,182,0,16,183,1,2,
/* out0407_em-eta7-phi20*/	7,62,1,3,62,2,4,73,0,4,73,1,3,74,0,2,74,2,3,182,1,16,
/* out0408_em-eta8-phi20*/	5,61,1,1,61,2,4,62,2,1,73,0,10,182,2,15,
/* out0409_em-eta9-phi20*/	8,61,0,1,61,2,10,72,0,2,8,1,4,8,2,2,50,0,5,50,2,4,182,2,1,
/* out0410_em-eta10-phi20*/	10,26,2,1,26,3,13,27,3,12,27,4,2,61,0,2,61,2,1,72,0,2,7,2,6,8,1,1,50,0,9,
/* out0411_em-eta11-phi20*/	9,26,0,2,26,1,5,26,2,15,26,3,3,27,0,7,27,4,5,7,1,10,7,2,3,49,0,1,
/* out0412_em-eta12-phi20*/	8,23,2,2,23,3,5,26,1,2,26,4,4,27,0,2,27,1,15,6,2,8,7,1,3,
/* out0413_em-eta13-phi20*/	8,22,2,1,23,2,4,23,3,9,23,4,11,23,5,1,6,0,4,6,1,3,6,2,3,
/* out0414_em-eta14-phi20*/	7,22,2,1,22,5,2,23,0,13,23,4,5,5,2,2,6,0,2,6,1,4,
/* out0415_em-eta15-phi20*/	7,10,3,1,22,4,13,22,5,1,23,1,3,1,1,1,5,0,5,5,2,1,
/* out0416_em-eta16-phi20*/	5,10,3,6,11,3,8,13,1,1,0,1,1,5,0,5,
/* out0417_em-eta17-phi20*/	5,11,2,2,11,3,7,11,4,3,0,1,5,5,0,1,
/* out0418_em-eta18-phi20*/	3,11,2,5,11,4,1,11,5,5,
/* out0419_em-eta19-phi20*/	2,8,4,4,11,5,5,
/* out0420_em-eta0-phi21*/	1,185,3,7,
/* out0421_em-eta1-phi21*/	2,185,2,9,185,3,9,
/* out0422_em-eta2-phi21*/	4,87,0,4,129,1,1,184,3,11,185,2,7,
/* out0423_em-eta3-phi21*/	8,86,1,6,86,2,4,87,0,5,87,1,14,129,0,12,129,1,2,184,2,12,184,3,5,
/* out0424_em-eta4-phi21*/	7,75,1,1,85,1,4,86,0,14,86,1,5,86,2,11,183,3,13,184,2,4,
/* out0425_em-eta5-phi21*/	7,74,1,1,75,2,2,85,0,15,85,1,6,85,2,3,183,2,14,183,3,3,
/* out0426_em-eta6-phi21*/	8,74,1,5,74,2,8,84,0,6,84,1,2,85,0,1,85,2,2,182,5,16,183,2,2,
/* out0427_em-eta7-phi21*/	5,73,1,12,73,2,1,74,2,2,84,0,4,182,4,16,
/* out0428_em-eta8-phi21*/	5,72,1,1,73,0,2,73,2,13,8,2,5,182,3,15,
/* out0429_em-eta9-phi21*/	6,72,0,5,72,1,8,8,0,6,8,1,5,8,2,9,182,3,1,
/* out0430_em-eta10-phi21*/	8,26,0,2,72,0,7,72,2,4,3,1,1,7,0,2,7,2,6,8,0,2,8,1,6,
/* out0431_em-eta11-phi21*/	7,25,2,13,25,5,5,26,0,12,26,1,4,7,0,11,7,1,1,7,2,1,
/* out0432_em-eta12-phi21*/	12,22,3,3,23,3,2,24,5,10,25,5,10,26,1,5,27,1,1,2,1,2,2,2,3,6,0,2,6,2,1,7,0,2,7,1,2,
/* out0433_em-eta13-phi21*/	7,22,0,6,22,2,6,22,3,13,24,5,1,1,2,1,2,1,2,6,0,7,
/* out0434_em-eta14-phi21*/	7,22,0,1,22,1,9,22,2,8,23,0,3,23,1,1,1,2,6,6,0,1,
/* out0435_em-eta15-phi21*/	5,10,0,4,10,3,1,22,1,1,23,1,11,1,1,6,
/* out0436_em-eta16-phi21*/	7,10,0,2,10,2,5,10,3,8,0,1,1,0,2,2,1,1,3,5,0,1,
/* out0437_em-eta17-phi21*/	5,10,2,5,11,0,1,11,4,7,0,1,5,0,2,1,
/* out0438_em-eta18-phi21*/	5,10,5,1,11,0,3,11,4,5,11,5,2,0,1,1,
/* out0439_em-eta19-phi21*/	2,10,5,6,11,5,4,
/* out0440_em-eta0-phi22*/	1,189,0,7,
/* out0441_em-eta1-phi22*/	2,189,0,9,189,1,9,
/* out0442_em-eta2-phi22*/	3,129,1,3,188,0,11,189,1,7,
/* out0443_em-eta3-phi22*/	8,127,1,4,128,1,1,128,2,6,129,0,4,129,1,10,129,2,16,188,0,5,188,1,12,
/* out0444_em-eta4-phi22*/	7,85,1,1,86,2,1,127,0,15,127,1,10,127,2,7,187,0,13,188,1,4,
/* out0445_em-eta5-phi22*/	8,85,1,5,85,2,10,126,0,9,126,1,3,127,0,1,127,2,1,187,0,3,187,1,14,
/* out0446_em-eta6-phi22*/	7,84,0,2,84,1,14,84,2,4,85,2,1,126,0,2,186,0,16,187,1,2,
/* out0447_em-eta7-phi22*/	7,73,1,1,73,2,1,83,0,1,83,1,5,84,0,4,84,2,9,186,1,16,
/* out0448_em-eta8-phi22*/	6,72,1,1,73,2,1,83,0,13,83,1,1,4,0,1,186,2,15,
/* out0449_em-eta9-phi22*/	8,72,1,6,72,2,4,83,0,2,3,2,3,4,0,2,4,1,12,8,0,7,186,2,1,
/* out0450_em-eta10-phi22*/	6,24,3,2,25,3,4,72,2,8,3,1,5,3,2,10,8,0,1,
/* out0451_em-eta11-phi22*/	9,24,2,6,24,3,4,25,2,3,25,3,12,25,4,12,25,5,1,2,2,5,3,1,8,7,0,1,
/* out0452_em-eta12-phi22*/	9,24,2,2,24,4,2,24,5,5,25,0,15,25,1,3,25,4,4,2,0,2,2,1,3,2,2,7,
/* out0453_em-eta13-phi22*/	4,22,0,6,24,4,13,1,2,1,2,1,8,
/* out0454_em-eta14-phi22*/	4,22,0,3,22,1,4,1,0,1,1,2,7,
/* out0455_em-eta15-phi22*/	6,10,0,5,22,1,2,23,1,1,1,0,3,1,1,3,1,2,1,
/* out0456_em-eta16-phi22*/	6,10,0,5,10,1,8,10,2,2,0,2,2,1,0,1,1,1,3,
/* out0457_em-eta17-phi22*/	5,10,1,1,10,2,4,11,0,6,11,1,1,0,2,6,
/* out0458_em-eta18-phi22*/	5,10,4,1,10,5,3,11,0,6,11,1,1,0,1,2,
/* out0459_em-eta19-phi22*/	2,10,4,2,10,5,6,
/* out0460_em-eta0-phi23*/	1,189,3,7,
/* out0461_em-eta1-phi23*/	2,189,2,9,189,3,9,
/* out0462_em-eta2-phi23*/	3,128,2,1,188,3,11,189,2,7,
/* out0463_em-eta3-phi23*/	5,128,0,16,128,1,13,128,2,9,188,2,12,188,3,5,
/* out0464_em-eta4-phi23*/	6,126,1,1,127,1,2,127,2,8,128,1,2,187,3,13,188,2,4,
/* out0465_em-eta5-phi23*/	5,126,0,3,126,1,12,126,2,11,187,2,14,187,3,3,
/* out0466_em-eta6-phi23*/	5,84,2,2,126,0,2,126,2,5,186,5,16,187,2,2,
/* out0467_em-eta7-phi23*/	3,83,1,7,84,2,1,186,4,16,
/* out0468_em-eta8-phi23*/	3,83,1,3,83,2,13,186,3,15,
/* out0469_em-eta9-phi23*/	5,83,2,3,3,2,1,4,0,13,4,1,4,186,3,1,
/* out0470_em-eta10-phi23*/	3,24,3,1,3,0,12,3,2,2,
/* out0471_em-eta11-phi23*/	8,24,0,15,24,1,2,24,2,4,24,3,9,2,0,1,2,2,1,3,0,4,3,1,2,
/* out0472_em-eta12-phi23*/	6,24,0,1,24,1,14,24,2,4,25,0,1,25,1,9,2,0,9,
/* out0473_em-eta13-phi23*/	4,24,4,1,25,1,4,2,0,4,2,1,1,
/* out0474_em-eta14-phi23*/	1,1,0,4,
/* out0475_em-eta15-phi23*/	1,1,0,6,
/* out0476_em-eta16-phi23*/	3,10,1,7,11,1,1,1,0,1,
/* out0477_em-eta17-phi23*/	2,11,1,11,0,2,3,
/* out0478_em-eta18-phi23*/	4,10,4,9,11,1,2,0,1,1,0,2,2,
/* out0479_em-eta19-phi23*/	1,10,4,4
};