parameter integer matrixH [0:5553] = {
/* num inputs = 180(in0-in179) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1691 */

/* out0000_had-eta0-phi0*/	1, 135, 0, 3, 
/* out0001_had-eta1-phi0*/	1, 135, 0, 4, 
/* out0002_had-eta2-phi0*/	2, 134, 0, 4, 135, 0, 1, 
/* out0003_had-eta3-phi0*/	1, 134, 0, 4, 
/* out0004_had-eta4-phi0*/	1, 133, 0, 4, 
/* out0005_had-eta5-phi0*/	5, 87, 0, 12, 87, 1, 4, 87, 2, 16, 94, 1, 2, 133, 0, 4, 
/* out0006_had-eta6-phi0*/	7, 86, 0, 5, 86, 2, 11, 87, 0, 2, 87, 1, 12, 93, 1, 1, 93, 2, 1, 132, 0, 3, 
/* out0007_had-eta7-phi0*/	5, 85, 2, 3, 86, 0, 6, 86, 1, 16, 86, 2, 5, 132, 0, 3, 
/* out0008_had-eta8-phi0*/	4, 85, 0, 6, 85, 1, 4, 85, 2, 13, 132, 0, 2, 
/* out0009_had-eta9-phi0*/	3, 84, 2, 7, 85, 0, 1, 85, 1, 9, 
/* out0010_had-eta10-phi0*/	3, 84, 0, 3, 84, 1, 5, 84, 2, 6, 
/* out0011_had-eta11-phi0*/	3, 83, 2, 5, 84, 1, 10, 127, 1, 5, 
/* out0012_had-eta12-phi0*/	5, 83, 0, 1, 83, 1, 2, 83, 2, 7, 126, 2, 2, 127, 1, 5, 
/* out0013_had-eta13-phi0*/	3, 83, 1, 8, 126, 1, 3, 126, 2, 6, 
/* out0014_had-eta14-phi0*/	3, 82, 2, 7, 83, 1, 1, 126, 1, 4, 
/* out0015_had-eta15-phi0*/	3, 82, 1, 3, 82, 2, 4, 125, 2, 5, 
/* out0016_had-eta16-phi0*/	3, 82, 1, 5, 125, 1, 4, 125, 2, 1, 
/* out0017_had-eta17-phi0*/	3, 81, 1, 3, 82, 1, 2, 125, 1, 1, 
/* out0018_had-eta18-phi0*/	2, 81, 1, 4, 124, 1, 2, 
/* out0019_had-eta19-phi0*/	2, 81, 1, 1, 124, 1, 2, 
/* out0020_had-eta0-phi1*/	1, 135, 0, 3, 
/* out0021_had-eta1-phi1*/	1, 135, 0, 4, 
/* out0022_had-eta2-phi1*/	2, 134, 0, 4, 135, 0, 1, 
/* out0023_had-eta3-phi1*/	1, 134, 0, 4, 
/* out0024_had-eta4-phi1*/	1, 133, 0, 4, 
/* out0025_had-eta5-phi1*/	6, 87, 0, 2, 93, 0, 2, 93, 2, 8, 94, 0, 13, 94, 1, 14, 133, 0, 4, 
/* out0026_had-eta6-phi1*/	5, 86, 0, 2, 93, 0, 5, 93, 1, 15, 93, 2, 7, 132, 0, 3, 
/* out0027_had-eta7-phi1*/	5, 86, 0, 3, 92, 0, 1, 92, 1, 5, 92, 2, 15, 132, 0, 3, 
/* out0028_had-eta8-phi1*/	4, 85, 0, 7, 91, 2, 5, 92, 1, 8, 132, 0, 2, 
/* out0029_had-eta9-phi1*/	6, 84, 0, 2, 84, 2, 3, 85, 0, 2, 85, 1, 3, 91, 1, 6, 91, 2, 6, 
/* out0030_had-eta10-phi1*/	3, 84, 0, 9, 90, 2, 2, 91, 1, 2, 
/* out0031_had-eta11-phi1*/	8, 83, 0, 1, 83, 2, 3, 84, 0, 2, 84, 1, 1, 90, 1, 3, 90, 2, 3, 127, 0, 10, 127, 1, 1, 
/* out0032_had-eta12-phi1*/	8, 83, 0, 9, 83, 2, 1, 90, 1, 1, 122, 2, 1, 126, 0, 2, 126, 2, 4, 127, 0, 5, 127, 1, 5, 
/* out0033_had-eta13-phi1*/	7, 82, 2, 1, 83, 0, 4, 83, 1, 3, 89, 2, 1, 126, 0, 6, 126, 1, 2, 126, 2, 4, 
/* out0034_had-eta14-phi1*/	6, 82, 0, 3, 82, 2, 3, 83, 1, 2, 125, 2, 2, 126, 0, 1, 126, 1, 7, 
/* out0035_had-eta15-phi1*/	5, 82, 0, 5, 82, 1, 1, 82, 2, 1, 125, 0, 1, 125, 2, 7, 
/* out0036_had-eta16-phi1*/	5, 82, 0, 1, 82, 1, 3, 125, 0, 1, 125, 1, 5, 125, 2, 1, 
/* out0037_had-eta17-phi1*/	4, 81, 1, 3, 82, 1, 1, 124, 1, 2, 125, 1, 4, 
/* out0038_had-eta18-phi1*/	3, 81, 0, 2, 81, 1, 3, 124, 1, 5, 
/* out0039_had-eta19-phi1*/	3, 81, 0, 1, 81, 1, 1, 124, 1, 1, 
/* out0040_had-eta0-phi2*/	1, 139, 0, 3, 
/* out0041_had-eta1-phi2*/	1, 139, 0, 4, 
/* out0042_had-eta2-phi2*/	2, 138, 0, 4, 139, 0, 1, 
/* out0043_had-eta3-phi2*/	1, 138, 0, 4, 
/* out0044_had-eta4-phi2*/	3, 70, 2, 1, 94, 0, 1, 137, 0, 4, 
/* out0045_had-eta5-phi2*/	6, 70, 0, 6, 70, 1, 13, 70, 2, 15, 93, 0, 1, 94, 0, 2, 137, 0, 4, 
/* out0046_had-eta6-phi2*/	5, 69, 1, 4, 69, 2, 14, 70, 1, 2, 93, 0, 8, 136, 0, 3, 
/* out0047_had-eta7-phi2*/	5, 68, 2, 3, 69, 1, 6, 92, 0, 13, 92, 2, 1, 136, 0, 3, 
/* out0048_had-eta8-phi2*/	7, 68, 1, 3, 68, 2, 3, 91, 0, 4, 91, 2, 4, 92, 0, 2, 92, 1, 3, 136, 0, 2, 
/* out0049_had-eta9-phi2*/	3, 91, 0, 10, 91, 1, 5, 91, 2, 1, 
/* out0050_had-eta10-phi2*/	3, 90, 0, 2, 90, 2, 8, 91, 1, 3, 
/* out0051_had-eta11-phi2*/	5, 90, 0, 2, 90, 1, 6, 90, 2, 3, 122, 2, 9, 127, 0, 1, 
/* out0052_had-eta12-phi2*/	5, 83, 0, 1, 89, 2, 4, 90, 1, 5, 122, 1, 8, 122, 2, 5, 
/* out0053_had-eta13-phi2*/	5, 89, 1, 1, 89, 2, 6, 121, 2, 3, 122, 1, 3, 126, 0, 5, 
/* out0054_had-eta14-phi2*/	5, 82, 0, 1, 89, 1, 6, 121, 1, 3, 121, 2, 4, 126, 0, 2, 
/* out0055_had-eta15-phi2*/	5, 82, 0, 4, 88, 2, 1, 89, 1, 1, 121, 1, 1, 125, 0, 7, 
/* out0056_had-eta16-phi2*/	3, 82, 0, 2, 88, 2, 3, 125, 0, 6, 
/* out0057_had-eta17-phi2*/	9, 81, 0, 4, 81, 1, 1, 82, 1, 1, 88, 1, 2, 120, 2, 1, 124, 0, 2, 124, 1, 2, 125, 0, 1, 125, 1, 2, 
/* out0058_had-eta18-phi2*/	3, 81, 0, 6, 124, 0, 5, 124, 1, 2, 
/* out0059_had-eta19-phi2*/	2, 81, 0, 1, 124, 0, 1, 
/* out0060_had-eta0-phi3*/	1, 139, 0, 3, 
/* out0061_had-eta1-phi3*/	1, 139, 0, 4, 
/* out0062_had-eta2-phi3*/	2, 138, 0, 4, 139, 0, 1, 
/* out0063_had-eta3-phi3*/	1, 138, 0, 4, 
/* out0064_had-eta4-phi3*/	1, 137, 0, 4, 
/* out0065_had-eta5-phi3*/	5, 70, 0, 10, 70, 1, 1, 73, 1, 3, 73, 2, 15, 137, 0, 4, 
/* out0066_had-eta6-phi3*/	6, 69, 0, 15, 69, 1, 1, 69, 2, 2, 72, 2, 3, 73, 1, 7, 136, 0, 3, 
/* out0067_had-eta7-phi3*/	7, 68, 0, 6, 68, 2, 8, 69, 0, 1, 69, 1, 5, 72, 1, 2, 72, 2, 2, 136, 0, 3, 
/* out0068_had-eta8-phi3*/	4, 68, 0, 4, 68, 1, 12, 68, 2, 2, 136, 0, 2, 
/* out0069_had-eta9-phi3*/	4, 67, 1, 1, 67, 2, 13, 68, 1, 1, 91, 0, 2, 
/* out0070_had-eta10-phi3*/	3, 67, 1, 8, 67, 2, 1, 90, 0, 4, 
/* out0071_had-eta11-phi3*/	4, 66, 2, 3, 90, 0, 8, 122, 0, 6, 122, 2, 1, 
/* out0072_had-eta12-phi3*/	8, 66, 1, 1, 66, 2, 1, 89, 0, 3, 89, 2, 3, 90, 1, 1, 122, 0, 10, 122, 1, 3, 123, 2, 1, 
/* out0073_had-eta13-phi3*/	6, 89, 0, 5, 89, 1, 1, 89, 2, 2, 121, 0, 3, 121, 2, 6, 122, 1, 2, 
/* out0074_had-eta14-phi3*/	4, 89, 1, 6, 121, 0, 2, 121, 1, 5, 121, 2, 3, 
/* out0075_had-eta15-phi3*/	3, 88, 2, 5, 120, 2, 2, 121, 1, 5, 
/* out0076_had-eta16-phi3*/	3, 88, 1, 1, 88, 2, 4, 120, 2, 6, 
/* out0077_had-eta17-phi3*/	4, 88, 1, 4, 120, 1, 4, 120, 2, 1, 124, 0, 1, 
/* out0078_had-eta18-phi3*/	4, 81, 0, 2, 88, 1, 1, 120, 1, 1, 124, 0, 7, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	1, 143, 0, 3, 
/* out0081_had-eta1-phi4*/	1, 143, 0, 4, 
/* out0082_had-eta2-phi4*/	2, 142, 0, 4, 143, 0, 1, 
/* out0083_had-eta3-phi4*/	1, 142, 0, 4, 
/* out0084_had-eta4-phi4*/	1, 141, 0, 4, 
/* out0085_had-eta5-phi4*/	5, 73, 0, 15, 73, 1, 1, 73, 2, 1, 74, 2, 7, 141, 0, 4, 
/* out0086_had-eta6-phi4*/	7, 72, 0, 8, 72, 2, 10, 73, 0, 1, 73, 1, 5, 74, 1, 3, 74, 2, 1, 140, 0, 3, 
/* out0087_had-eta7-phi4*/	6, 68, 0, 2, 71, 2, 4, 72, 0, 3, 72, 1, 14, 72, 2, 1, 140, 0, 3, 
/* out0088_had-eta8-phi4*/	5, 67, 2, 1, 68, 0, 4, 71, 1, 5, 71, 2, 9, 140, 0, 2, 
/* out0089_had-eta9-phi4*/	3, 67, 0, 13, 67, 2, 1, 71, 1, 2, 
/* out0090_had-eta10-phi4*/	4, 66, 0, 1, 66, 2, 3, 67, 0, 3, 67, 1, 7, 
/* out0091_had-eta11-phi4*/	4, 66, 0, 1, 66, 1, 1, 66, 2, 9, 123, 2, 4, 
/* out0092_had-eta12-phi4*/	4, 66, 1, 9, 89, 0, 1, 123, 1, 2, 123, 2, 11, 
/* out0093_had-eta13-phi4*/	4, 60, 2, 2, 89, 0, 5, 121, 0, 4, 123, 1, 7, 
/* out0094_had-eta14-phi4*/	6, 60, 1, 1, 60, 2, 2, 89, 0, 2, 89, 1, 1, 116, 2, 2, 121, 0, 7, 
/* out0095_had-eta15-phi4*/	6, 88, 0, 4, 88, 2, 2, 116, 2, 1, 120, 0, 2, 120, 2, 3, 121, 1, 2, 
/* out0096_had-eta16-phi4*/	5, 88, 0, 3, 88, 1, 1, 88, 2, 1, 120, 0, 3, 120, 2, 3, 
/* out0097_had-eta17-phi4*/	2, 88, 1, 4, 120, 1, 5, 
/* out0098_had-eta18-phi4*/	2, 88, 1, 1, 120, 1, 3, 
/* out0099_had-eta19-phi4*/	0, 
/* out0100_had-eta0-phi5*/	1, 143, 0, 3, 
/* out0101_had-eta1-phi5*/	1, 143, 0, 4, 
/* out0102_had-eta2-phi5*/	2, 142, 0, 4, 143, 0, 1, 
/* out0103_had-eta3-phi5*/	1, 142, 0, 4, 
/* out0104_had-eta4-phi5*/	1, 141, 0, 4, 
/* out0105_had-eta5-phi5*/	4, 74, 0, 14, 74, 1, 1, 74, 2, 8, 141, 0, 4, 
/* out0106_had-eta6-phi5*/	5, 72, 0, 3, 74, 0, 2, 74, 1, 12, 77, 2, 10, 140, 0, 3, 
/* out0107_had-eta7-phi5*/	6, 71, 0, 5, 71, 2, 2, 72, 0, 2, 77, 1, 8, 77, 2, 6, 140, 0, 3, 
/* out0108_had-eta8-phi5*/	4, 71, 0, 11, 71, 1, 6, 71, 2, 1, 140, 0, 2, 
/* out0109_had-eta9-phi5*/	2, 71, 1, 3, 75, 2, 12, 
/* out0110_had-eta10-phi5*/	3, 66, 0, 2, 75, 1, 8, 75, 2, 4, 
/* out0111_had-eta11-phi5*/	2, 66, 0, 10, 123, 0, 3, 
/* out0112_had-eta12-phi5*/	5, 60, 2, 2, 66, 0, 2, 66, 1, 5, 123, 0, 12, 123, 1, 1, 
/* out0113_had-eta13-phi5*/	4, 60, 2, 8, 116, 2, 5, 123, 0, 1, 123, 1, 6, 
/* out0114_had-eta14-phi5*/	4, 60, 1, 5, 60, 2, 2, 116, 1, 1, 116, 2, 8, 
/* out0115_had-eta15-phi5*/	4, 60, 1, 2, 88, 0, 3, 116, 1, 6, 120, 0, 2, 
/* out0116_had-eta16-phi5*/	2, 88, 0, 4, 120, 0, 6, 
/* out0117_had-eta17-phi5*/	4, 88, 0, 2, 88, 1, 2, 120, 0, 3, 120, 1, 2, 
/* out0118_had-eta18-phi5*/	1, 120, 1, 1, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	1, 147, 0, 3, 
/* out0121_had-eta1-phi6*/	1, 147, 0, 4, 
/* out0122_had-eta2-phi6*/	2, 146, 0, 4, 147, 0, 1, 
/* out0123_had-eta3-phi6*/	1, 146, 0, 4, 
/* out0124_had-eta4-phi6*/	1, 145, 0, 4, 
/* out0125_had-eta5-phi6*/	4, 79, 0, 8, 79, 1, 1, 79, 2, 14, 145, 0, 4, 
/* out0126_had-eta6-phi6*/	5, 77, 0, 10, 78, 2, 3, 79, 1, 12, 79, 2, 2, 144, 0, 3, 
/* out0127_had-eta7-phi6*/	6, 76, 0, 2, 76, 2, 5, 77, 0, 6, 77, 1, 8, 78, 2, 2, 144, 0, 3, 
/* out0128_had-eta8-phi6*/	4, 76, 0, 1, 76, 1, 6, 76, 2, 11, 144, 0, 2, 
/* out0129_had-eta9-phi6*/	2, 75, 0, 12, 76, 1, 3, 
/* out0130_had-eta10-phi6*/	3, 61, 2, 2, 75, 0, 4, 75, 1, 8, 
/* out0131_had-eta11-phi6*/	2, 61, 2, 10, 118, 2, 3, 
/* out0132_had-eta12-phi6*/	5, 60, 0, 2, 61, 1, 5, 61, 2, 2, 118, 1, 1, 118, 2, 12, 
/* out0133_had-eta13-phi6*/	4, 60, 0, 7, 116, 0, 5, 118, 1, 6, 118, 2, 1, 
/* out0134_had-eta14-phi6*/	4, 60, 0, 2, 60, 1, 5, 116, 0, 8, 116, 1, 1, 
/* out0135_had-eta15-phi6*/	4, 53, 2, 3, 60, 1, 2, 115, 2, 2, 116, 1, 7, 
/* out0136_had-eta16-phi6*/	2, 53, 2, 4, 115, 2, 6, 
/* out0137_had-eta17-phi6*/	4, 53, 1, 2, 53, 2, 2, 115, 1, 2, 115, 2, 3, 
/* out0138_had-eta18-phi6*/	1, 115, 1, 1, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	1, 147, 0, 3, 
/* out0141_had-eta1-phi7*/	1, 147, 0, 4, 
/* out0142_had-eta2-phi7*/	2, 146, 0, 4, 147, 0, 1, 
/* out0143_had-eta3-phi7*/	1, 146, 0, 4, 
/* out0144_had-eta4-phi7*/	1, 145, 0, 4, 
/* out0145_had-eta5-phi7*/	5, 79, 0, 7, 80, 0, 1, 80, 1, 1, 80, 2, 15, 145, 0, 4, 
/* out0146_had-eta6-phi7*/	7, 78, 0, 10, 78, 2, 8, 79, 0, 1, 79, 1, 3, 80, 1, 5, 80, 2, 1, 144, 0, 3, 
/* out0147_had-eta7-phi7*/	6, 63, 2, 2, 76, 0, 4, 78, 0, 1, 78, 1, 14, 78, 2, 3, 144, 0, 3, 
/* out0148_had-eta8-phi7*/	5, 62, 0, 1, 63, 2, 4, 76, 0, 9, 76, 1, 5, 144, 0, 2, 
/* out0149_had-eta9-phi7*/	3, 62, 0, 1, 62, 2, 13, 76, 1, 2, 
/* out0150_had-eta10-phi7*/	4, 61, 0, 3, 61, 2, 1, 62, 1, 7, 62, 2, 3, 
/* out0151_had-eta11-phi7*/	4, 61, 0, 9, 61, 1, 1, 61, 2, 1, 118, 0, 4, 
/* out0152_had-eta12-phi7*/	4, 54, 2, 1, 61, 1, 9, 118, 0, 11, 118, 1, 2, 
/* out0153_had-eta13-phi7*/	4, 54, 2, 5, 60, 0, 3, 117, 2, 4, 118, 1, 7, 
/* out0154_had-eta14-phi7*/	7, 53, 0, 1, 54, 1, 1, 54, 2, 2, 60, 0, 2, 60, 1, 1, 116, 0, 2, 117, 2, 7, 
/* out0155_had-eta15-phi7*/	7, 53, 0, 2, 53, 2, 4, 115, 0, 3, 115, 2, 2, 116, 0, 1, 116, 1, 1, 117, 1, 2, 
/* out0156_had-eta16-phi7*/	5, 53, 0, 1, 53, 1, 1, 53, 2, 3, 115, 0, 3, 115, 2, 3, 
/* out0157_had-eta17-phi7*/	2, 53, 1, 4, 115, 1, 5, 
/* out0158_had-eta18-phi7*/	2, 53, 1, 1, 115, 1, 3, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	1, 151, 0, 3, 
/* out0161_had-eta1-phi8*/	1, 151, 0, 4, 
/* out0162_had-eta2-phi8*/	2, 150, 0, 4, 151, 0, 1, 
/* out0163_had-eta3-phi8*/	1, 150, 0, 4, 
/* out0164_had-eta4-phi8*/	1, 149, 0, 4, 
/* out0165_had-eta5-phi8*/	5, 65, 1, 1, 65, 2, 10, 80, 0, 15, 80, 1, 3, 149, 0, 4, 
/* out0166_had-eta6-phi8*/	6, 64, 0, 2, 64, 1, 1, 64, 2, 15, 78, 0, 3, 80, 1, 7, 148, 0, 3, 
/* out0167_had-eta7-phi8*/	7, 63, 0, 8, 63, 2, 6, 64, 1, 5, 64, 2, 1, 78, 0, 2, 78, 1, 2, 148, 0, 3, 
/* out0168_had-eta8-phi8*/	4, 63, 0, 2, 63, 1, 12, 63, 2, 4, 148, 0, 2, 
/* out0169_had-eta9-phi8*/	4, 56, 2, 2, 62, 0, 13, 62, 1, 1, 63, 1, 1, 
/* out0170_had-eta10-phi8*/	3, 55, 2, 4, 62, 0, 1, 62, 1, 8, 
/* out0171_had-eta11-phi8*/	4, 55, 2, 8, 61, 0, 3, 119, 0, 1, 119, 2, 6, 
/* out0172_had-eta12-phi8*/	8, 54, 0, 3, 54, 2, 3, 55, 1, 1, 61, 0, 1, 61, 1, 1, 118, 0, 1, 119, 1, 3, 119, 2, 10, 
/* out0173_had-eta13-phi8*/	6, 54, 0, 2, 54, 1, 1, 54, 2, 5, 117, 0, 6, 117, 2, 3, 119, 1, 2, 
/* out0174_had-eta14-phi8*/	4, 54, 1, 6, 117, 0, 3, 117, 1, 5, 117, 2, 2, 
/* out0175_had-eta15-phi8*/	3, 53, 0, 5, 115, 0, 2, 117, 1, 5, 
/* out0176_had-eta16-phi8*/	3, 53, 0, 3, 53, 1, 1, 115, 0, 6, 
/* out0177_had-eta17-phi8*/	4, 53, 1, 4, 111, 1, 1, 115, 0, 1, 115, 1, 4, 
/* out0178_had-eta18-phi8*/	4, 46, 1, 3, 53, 1, 1, 111, 1, 7, 115, 1, 1, 
/* out0179_had-eta19-phi8*/	0, 
/* out0180_had-eta0-phi9*/	1, 151, 0, 3, 
/* out0181_had-eta1-phi9*/	1, 151, 0, 4, 
/* out0182_had-eta2-phi9*/	2, 150, 0, 4, 151, 0, 1, 
/* out0183_had-eta3-phi9*/	1, 150, 0, 4, 
/* out0184_had-eta4-phi9*/	3, 59, 1, 1, 65, 0, 1, 149, 0, 4, 
/* out0185_had-eta5-phi9*/	6, 58, 2, 1, 59, 1, 2, 65, 0, 15, 65, 1, 13, 65, 2, 6, 149, 0, 4, 
/* out0186_had-eta6-phi9*/	5, 58, 2, 8, 64, 0, 14, 64, 1, 4, 65, 1, 2, 148, 0, 3, 
/* out0187_had-eta7-phi9*/	5, 57, 0, 1, 57, 2, 13, 63, 0, 3, 64, 1, 6, 148, 0, 3, 
/* out0188_had-eta8-phi9*/	7, 56, 0, 4, 56, 2, 4, 57, 1, 3, 57, 2, 2, 63, 0, 3, 63, 1, 3, 148, 0, 2, 
/* out0189_had-eta9-phi9*/	3, 56, 0, 1, 56, 1, 5, 56, 2, 10, 
/* out0190_had-eta10-phi9*/	3, 55, 0, 8, 55, 2, 2, 56, 1, 3, 
/* out0191_had-eta11-phi9*/	5, 55, 0, 3, 55, 1, 6, 55, 2, 2, 114, 1, 1, 119, 0, 9, 
/* out0192_had-eta12-phi9*/	5, 48, 2, 1, 54, 0, 4, 55, 1, 5, 119, 0, 5, 119, 1, 8, 
/* out0193_had-eta13-phi9*/	5, 54, 0, 6, 54, 1, 1, 113, 2, 5, 117, 0, 3, 119, 1, 3, 
/* out0194_had-eta14-phi9*/	5, 47, 2, 1, 54, 1, 6, 113, 2, 2, 117, 0, 4, 117, 1, 3, 
/* out0195_had-eta15-phi9*/	5, 47, 2, 4, 53, 0, 1, 54, 1, 1, 112, 2, 7, 117, 1, 1, 
/* out0196_had-eta16-phi9*/	3, 47, 2, 2, 53, 0, 3, 112, 2, 6, 
/* out0197_had-eta17-phi9*/	7, 46, 1, 4, 53, 1, 2, 111, 0, 2, 111, 1, 2, 112, 1, 2, 112, 2, 1, 115, 0, 1, 
/* out0198_had-eta18-phi9*/	3, 46, 1, 6, 111, 0, 2, 111, 1, 5, 
/* out0199_had-eta19-phi9*/	1, 111, 1, 1, 
/* out0200_had-eta0-phi10*/	1, 155, 0, 3, 
/* out0201_had-eta1-phi10*/	1, 155, 0, 4, 
/* out0202_had-eta2-phi10*/	2, 154, 0, 4, 155, 0, 1, 
/* out0203_had-eta3-phi10*/	1, 154, 0, 4, 
/* out0204_had-eta4-phi10*/	1, 153, 0, 4, 
/* out0205_had-eta5-phi10*/	6, 52, 2, 2, 58, 0, 8, 58, 2, 2, 59, 0, 14, 59, 1, 13, 153, 0, 4, 
/* out0206_had-eta6-phi10*/	5, 51, 2, 2, 58, 0, 7, 58, 1, 15, 58, 2, 5, 152, 0, 3, 
/* out0207_had-eta7-phi10*/	5, 51, 2, 3, 57, 0, 15, 57, 1, 5, 57, 2, 1, 152, 0, 3, 
/* out0208_had-eta8-phi10*/	4, 50, 2, 7, 56, 0, 5, 57, 1, 8, 152, 0, 2, 
/* out0209_had-eta9-phi10*/	4, 49, 2, 2, 50, 2, 2, 56, 0, 6, 56, 1, 6, 
/* out0210_had-eta10-phi10*/	3, 49, 2, 9, 55, 0, 2, 56, 1, 2, 
/* out0211_had-eta11-phi10*/	8, 48, 0, 1, 48, 2, 1, 49, 1, 1, 49, 2, 2, 55, 0, 3, 55, 1, 3, 114, 0, 1, 114, 1, 10, 
/* out0212_had-eta12-phi10*/	7, 48, 2, 9, 55, 1, 1, 113, 0, 4, 113, 2, 2, 114, 0, 5, 114, 1, 5, 119, 0, 1, 
/* out0213_had-eta13-phi10*/	6, 48, 1, 2, 48, 2, 4, 54, 0, 1, 113, 0, 4, 113, 1, 2, 113, 2, 6, 
/* out0214_had-eta14-phi10*/	5, 47, 0, 3, 47, 2, 3, 112, 0, 2, 113, 1, 7, 113, 2, 1, 
/* out0215_had-eta15-phi10*/	3, 47, 2, 5, 112, 0, 7, 112, 2, 1, 
/* out0216_had-eta16-phi10*/	5, 47, 1, 3, 47, 2, 1, 112, 0, 1, 112, 1, 5, 112, 2, 1, 
/* out0217_had-eta17-phi10*/	4, 46, 0, 3, 47, 1, 1, 111, 0, 2, 112, 1, 4, 
/* out0218_had-eta18-phi10*/	3, 46, 0, 2, 46, 1, 2, 111, 0, 5, 
/* out0219_had-eta19-phi10*/	2, 46, 1, 1, 111, 0, 1, 
/* out0220_had-eta0-phi11*/	1, 155, 0, 3, 
/* out0221_had-eta1-phi11*/	1, 155, 0, 4, 
/* out0222_had-eta2-phi11*/	2, 154, 0, 4, 155, 0, 1, 
/* out0223_had-eta3-phi11*/	1, 154, 0, 4, 
/* out0224_had-eta4-phi11*/	1, 153, 0, 4, 
/* out0225_had-eta5-phi11*/	5, 52, 0, 12, 52, 1, 4, 52, 2, 12, 59, 0, 2, 153, 0, 4, 
/* out0226_had-eta6-phi11*/	7, 51, 0, 11, 51, 2, 5, 52, 1, 8, 52, 2, 2, 58, 0, 1, 58, 1, 1, 152, 0, 3, 
/* out0227_had-eta7-phi11*/	5, 50, 0, 3, 51, 0, 1, 51, 1, 12, 51, 2, 6, 152, 0, 3, 
/* out0228_had-eta8-phi11*/	4, 50, 0, 9, 50, 1, 4, 50, 2, 6, 152, 0, 2, 
/* out0229_had-eta9-phi11*/	3, 49, 0, 7, 50, 1, 8, 50, 2, 1, 
/* out0230_had-eta10-phi11*/	3, 49, 0, 5, 49, 1, 5, 49, 2, 3, 
/* out0231_had-eta11-phi11*/	3, 48, 0, 5, 49, 1, 6, 114, 0, 5, 
/* out0232_had-eta12-phi11*/	6, 48, 0, 7, 48, 1, 2, 48, 2, 1, 110, 2, 6, 113, 0, 2, 114, 0, 5, 
/* out0233_had-eta13-phi11*/	4, 48, 1, 8, 110, 2, 2, 113, 0, 6, 113, 1, 3, 
/* out0234_had-eta14-phi11*/	4, 47, 0, 6, 48, 1, 1, 109, 2, 4, 113, 1, 4, 
/* out0235_had-eta15-phi11*/	4, 47, 0, 3, 47, 1, 2, 109, 2, 3, 112, 0, 5, 
/* out0236_had-eta16-phi11*/	4, 47, 1, 5, 108, 2, 1, 112, 0, 1, 112, 1, 4, 
/* out0237_had-eta17-phi11*/	4, 46, 0, 3, 47, 1, 1, 108, 2, 4, 112, 1, 1, 
/* out0238_had-eta18-phi11*/	3, 46, 0, 3, 108, 2, 3, 111, 0, 2, 
/* out0239_had-eta19-phi11*/	2, 46, 0, 1, 111, 0, 2, 
/* out0240_had-eta0-phi12*/	1, 159, 0, 3, 
/* out0241_had-eta1-phi12*/	1, 159, 0, 4, 
/* out0242_had-eta2-phi12*/	2, 158, 0, 4, 159, 0, 1, 
/* out0243_had-eta3-phi12*/	1, 158, 0, 4, 
/* out0244_had-eta4-phi12*/	1, 157, 0, 4, 
/* out0245_had-eta5-phi12*/	7, 44, 0, 5, 44, 2, 1, 45, 0, 9, 45, 1, 16, 52, 0, 4, 52, 1, 3, 157, 0, 4, 
/* out0246_had-eta6-phi12*/	6, 44, 0, 3, 44, 1, 6, 44, 2, 15, 51, 0, 3, 52, 1, 1, 156, 0, 3, 
/* out0247_had-eta7-phi12*/	6, 43, 0, 5, 43, 2, 11, 44, 1, 1, 51, 0, 1, 51, 1, 4, 156, 0, 3, 
/* out0248_had-eta8-phi12*/	7, 42, 0, 2, 42, 2, 1, 43, 1, 4, 43, 2, 5, 50, 0, 4, 50, 1, 2, 156, 0, 2, 
/* out0249_had-eta9-phi12*/	4, 42, 0, 1, 42, 2, 12, 49, 0, 1, 50, 1, 2, 
/* out0250_had-eta10-phi12*/	6, 41, 0, 1, 41, 2, 2, 42, 1, 2, 42, 2, 2, 49, 0, 3, 49, 1, 3, 
/* out0251_had-eta11-phi12*/	3, 41, 2, 9, 49, 1, 1, 110, 0, 5, 
/* out0252_had-eta12-phi12*/	7, 41, 1, 1, 41, 2, 3, 48, 0, 3, 48, 1, 1, 110, 0, 5, 110, 1, 2, 110, 2, 6, 
/* out0253_had-eta13-phi12*/	5, 40, 2, 5, 48, 1, 2, 109, 0, 3, 110, 1, 6, 110, 2, 2, 
/* out0254_had-eta14-phi12*/	4, 40, 2, 5, 47, 0, 2, 109, 0, 4, 109, 2, 5, 
/* out0255_had-eta15-phi12*/	5, 40, 2, 1, 47, 0, 2, 47, 1, 2, 109, 1, 5, 109, 2, 4, 
/* out0256_had-eta16-phi12*/	5, 39, 2, 3, 47, 1, 2, 108, 0, 4, 108, 2, 1, 109, 1, 1, 
/* out0257_had-eta17-phi12*/	4, 39, 2, 3, 46, 0, 1, 108, 0, 1, 108, 2, 4, 
/* out0258_had-eta18-phi12*/	4, 39, 2, 1, 46, 0, 2, 108, 1, 2, 108, 2, 3, 
/* out0259_had-eta19-phi12*/	2, 46, 0, 1, 108, 1, 2, 
/* out0260_had-eta0-phi13*/	1, 159, 0, 3, 
/* out0261_had-eta1-phi13*/	1, 159, 0, 4, 
/* out0262_had-eta2-phi13*/	2, 158, 0, 4, 159, 0, 1, 
/* out0263_had-eta3-phi13*/	1, 158, 0, 4, 
/* out0264_had-eta4-phi13*/	1, 157, 0, 4, 
/* out0265_had-eta5-phi13*/	6, 38, 0, 7, 38, 1, 2, 38, 2, 14, 44, 0, 3, 45, 0, 7, 157, 0, 4, 
/* out0266_had-eta6-phi13*/	7, 37, 0, 2, 37, 2, 7, 38, 1, 2, 38, 2, 2, 44, 0, 5, 44, 1, 9, 156, 0, 3, 
/* out0267_had-eta7-phi13*/	5, 36, 2, 1, 37, 2, 7, 43, 0, 11, 43, 1, 4, 156, 0, 3, 
/* out0268_had-eta8-phi13*/	4, 36, 2, 7, 42, 0, 5, 43, 1, 8, 156, 0, 2, 
/* out0269_had-eta9-phi13*/	3, 42, 0, 8, 42, 1, 8, 42, 2, 1, 
/* out0270_had-eta10-phi13*/	3, 35, 2, 1, 41, 0, 7, 42, 1, 5, 
/* out0271_had-eta11-phi13*/	5, 41, 0, 5, 41, 1, 4, 41, 2, 2, 107, 1, 10, 110, 0, 1, 
/* out0272_had-eta12-phi13*/	7, 40, 0, 3, 41, 1, 6, 105, 2, 2, 107, 0, 1, 107, 1, 5, 110, 0, 5, 110, 1, 4, 
/* out0273_had-eta13-phi13*/	5, 40, 0, 5, 40, 2, 2, 105, 2, 6, 109, 0, 2, 110, 1, 4, 
/* out0274_had-eta14-phi13*/	5, 40, 1, 4, 40, 2, 3, 105, 2, 1, 109, 0, 7, 109, 1, 2, 
/* out0275_had-eta15-phi13*/	4, 39, 0, 2, 40, 1, 3, 103, 2, 1, 109, 1, 7, 
/* out0276_had-eta16-phi13*/	5, 39, 0, 2, 39, 2, 3, 103, 2, 1, 108, 0, 5, 109, 1, 1, 
/* out0277_had-eta17-phi13*/	3, 39, 2, 4, 108, 0, 4, 108, 1, 2, 
/* out0278_had-eta18-phi13*/	3, 39, 1, 1, 39, 2, 2, 108, 1, 5, 
/* out0279_had-eta19-phi13*/	2, 39, 1, 1, 108, 1, 1, 
/* out0280_had-eta0-phi14*/	1, 163, 0, 3, 
/* out0281_had-eta1-phi14*/	1, 163, 0, 4, 
/* out0282_had-eta2-phi14*/	2, 162, 0, 4, 163, 0, 1, 
/* out0283_had-eta3-phi14*/	1, 162, 0, 4, 
/* out0284_had-eta4-phi14*/	1, 161, 0, 4, 
/* out0285_had-eta5-phi14*/	5, 32, 0, 2, 32, 2, 6, 38, 0, 9, 38, 1, 9, 161, 0, 4, 
/* out0286_had-eta6-phi14*/	6, 32, 2, 7, 37, 0, 14, 37, 1, 4, 37, 2, 1, 38, 1, 3, 160, 0, 3, 
/* out0287_had-eta7-phi14*/	5, 31, 2, 3, 36, 0, 8, 37, 1, 12, 37, 2, 1, 160, 0, 3, 
/* out0288_had-eta8-phi14*/	4, 36, 0, 5, 36, 1, 7, 36, 2, 7, 160, 0, 2, 
/* out0289_had-eta9-phi14*/	5, 35, 0, 6, 35, 2, 4, 36, 1, 3, 36, 2, 1, 42, 1, 1, 
/* out0290_had-eta10-phi14*/	3, 35, 1, 2, 35, 2, 10, 41, 0, 1, 
/* out0291_had-eta11-phi14*/	8, 34, 0, 1, 34, 2, 3, 35, 1, 1, 35, 2, 1, 41, 0, 2, 41, 1, 3, 107, 0, 9, 107, 1, 1, 
/* out0292_had-eta12-phi14*/	5, 34, 2, 6, 40, 0, 2, 41, 1, 2, 105, 0, 8, 107, 0, 5, 
/* out0293_had-eta13-phi14*/	6, 34, 2, 1, 40, 0, 6, 40, 1, 1, 105, 0, 3, 105, 1, 3, 105, 2, 5, 
/* out0294_had-eta14-phi14*/	4, 40, 1, 6, 103, 0, 3, 105, 1, 4, 105, 2, 2, 
/* out0295_had-eta15-phi14*/	4, 39, 0, 4, 40, 1, 2, 103, 0, 1, 103, 2, 7, 
/* out0296_had-eta16-phi14*/	2, 39, 0, 4, 103, 2, 6, 
/* out0297_had-eta17-phi14*/	6, 39, 1, 4, 102, 2, 1, 103, 1, 1, 103, 2, 1, 108, 0, 2, 108, 1, 2, 
/* out0298_had-eta18-phi14*/	3, 39, 1, 3, 102, 2, 4, 108, 1, 2, 
/* out0299_had-eta19-phi14*/	1, 102, 2, 2, 
/* out0300_had-eta0-phi15*/	1, 163, 0, 3, 
/* out0301_had-eta1-phi15*/	1, 163, 0, 4, 
/* out0302_had-eta2-phi15*/	2, 162, 0, 4, 163, 0, 1, 
/* out0303_had-eta3-phi15*/	1, 162, 0, 4, 
/* out0304_had-eta4-phi15*/	2, 28, 1, 1, 161, 0, 4, 
/* out0305_had-eta5-phi15*/	6, 26, 2, 1, 28, 1, 14, 32, 0, 14, 32, 1, 3, 32, 2, 1, 161, 0, 4, 
/* out0306_had-eta6-phi15*/	6, 26, 2, 2, 31, 0, 10, 31, 2, 1, 32, 1, 13, 32, 2, 2, 160, 0, 3, 
/* out0307_had-eta7-phi15*/	5, 31, 0, 3, 31, 1, 7, 31, 2, 12, 36, 0, 1, 160, 0, 3, 
/* out0308_had-eta8-phi15*/	6, 30, 0, 4, 30, 2, 8, 31, 1, 1, 36, 0, 2, 36, 1, 5, 160, 0, 2, 
/* out0309_had-eta9-phi15*/	4, 30, 2, 6, 35, 0, 9, 35, 1, 1, 36, 1, 1, 
/* out0310_had-eta10-phi15*/	3, 29, 2, 1, 35, 0, 1, 35, 1, 11, 
/* out0311_had-eta11-phi15*/	6, 34, 0, 10, 34, 2, 1, 35, 1, 1, 106, 0, 7, 106, 2, 6, 107, 0, 1, 
/* out0312_had-eta12-phi15*/	6, 34, 0, 1, 34, 1, 4, 34, 2, 4, 105, 0, 3, 106, 1, 1, 106, 2, 10, 
/* out0313_had-eta13-phi15*/	7, 33, 0, 2, 33, 2, 1, 34, 1, 3, 34, 2, 1, 104, 2, 3, 105, 0, 2, 105, 1, 6, 
/* out0314_had-eta14-phi15*/	4, 33, 2, 6, 103, 0, 5, 104, 2, 2, 105, 1, 3, 
/* out0315_had-eta15-phi15*/	4, 33, 2, 5, 39, 0, 1, 103, 0, 5, 103, 1, 2, 
/* out0316_had-eta16-phi15*/	3, 39, 0, 3, 39, 1, 1, 103, 1, 6, 
/* out0317_had-eta17-phi15*/	4, 39, 1, 4, 102, 0, 4, 102, 2, 1, 103, 1, 1, 
/* out0318_had-eta18-phi15*/	3, 39, 1, 2, 102, 0, 1, 102, 2, 5, 
/* out0319_had-eta19-phi15*/	1, 102, 2, 3, 
/* out0320_had-eta0-phi16*/	1, 167, 0, 3, 
/* out0321_had-eta1-phi16*/	1, 167, 0, 4, 
/* out0322_had-eta2-phi16*/	2, 166, 0, 4, 167, 0, 1, 
/* out0323_had-eta3-phi16*/	1, 166, 0, 4, 
/* out0324_had-eta4-phi16*/	1, 165, 0, 4, 
/* out0325_had-eta5-phi16*/	6, 26, 0, 12, 26, 2, 1, 27, 1, 7, 28, 0, 16, 28, 1, 1, 165, 0, 4, 
/* out0326_had-eta6-phi16*/	6, 25, 0, 1, 26, 0, 2, 26, 1, 10, 26, 2, 12, 31, 0, 2, 164, 0, 3, 
/* out0327_had-eta7-phi16*/	6, 25, 0, 3, 25, 2, 11, 30, 0, 1, 31, 0, 1, 31, 1, 8, 164, 0, 3, 
/* out0328_had-eta8-phi16*/	5, 25, 2, 2, 30, 0, 11, 30, 1, 5, 30, 2, 1, 164, 0, 2, 
/* out0329_had-eta9-phi16*/	3, 29, 0, 5, 30, 1, 9, 30, 2, 1, 
/* out0330_had-eta10-phi16*/	2, 29, 0, 3, 29, 2, 10, 
/* out0331_had-eta11-phi16*/	6, 29, 1, 1, 29, 2, 5, 34, 0, 4, 34, 1, 1, 106, 0, 9, 106, 1, 4, 
/* out0332_had-eta12-phi16*/	4, 14, 2, 2, 34, 1, 7, 104, 0, 2, 106, 1, 11, 
/* out0333_had-eta13-phi16*/	5, 14, 2, 1, 33, 0, 6, 34, 1, 1, 104, 0, 7, 104, 2, 4, 
/* out0334_had-eta14-phi16*/	5, 33, 0, 4, 33, 1, 1, 33, 2, 1, 104, 1, 2, 104, 2, 7, 
/* out0335_had-eta15-phi16*/	6, 33, 1, 4, 33, 2, 2, 98, 2, 1, 103, 0, 2, 103, 1, 3, 104, 1, 1, 
/* out0336_had-eta16-phi16*/	6, 0, 0, 1, 0, 2, 1, 33, 1, 1, 33, 2, 1, 98, 2, 3, 103, 1, 3, 
/* out0337_had-eta17-phi16*/	2, 0, 2, 4, 102, 0, 5, 
/* out0338_had-eta18-phi16*/	3, 0, 2, 4, 102, 0, 3, 102, 1, 2, 
/* out0339_had-eta19-phi16*/	1, 102, 1, 4, 
/* out0340_had-eta0-phi17*/	1, 167, 0, 3, 
/* out0341_had-eta1-phi17*/	1, 167, 0, 4, 
/* out0342_had-eta2-phi17*/	2, 166, 0, 4, 167, 0, 1, 
/* out0343_had-eta3-phi17*/	1, 166, 0, 4, 
/* out0344_had-eta4-phi17*/	1, 165, 0, 4, 
/* out0345_had-eta5-phi17*/	5, 23, 0, 5, 26, 0, 2, 27, 0, 16, 27, 1, 9, 165, 0, 4, 
/* out0346_had-eta6-phi17*/	5, 23, 0, 2, 23, 2, 15, 25, 0, 4, 26, 1, 6, 164, 0, 3, 
/* out0347_had-eta7-phi17*/	4, 25, 0, 8, 25, 1, 13, 25, 2, 2, 164, 0, 3, 
/* out0348_had-eta8-phi17*/	6, 19, 0, 8, 19, 2, 5, 25, 1, 3, 25, 2, 1, 30, 1, 1, 164, 0, 2, 
/* out0349_had-eta9-phi17*/	3, 19, 2, 11, 29, 0, 5, 30, 1, 1, 
/* out0350_had-eta10-phi17*/	2, 29, 0, 3, 29, 1, 10, 
/* out0351_had-eta11-phi17*/	4, 14, 0, 6, 29, 1, 5, 101, 0, 7, 101, 2, 3, 
/* out0352_had-eta12-phi17*/	4, 14, 0, 2, 14, 2, 8, 101, 2, 12, 104, 0, 1, 
/* out0353_had-eta13-phi17*/	5, 14, 2, 5, 33, 0, 2, 101, 2, 1, 104, 0, 6, 104, 1, 5, 
/* out0354_had-eta14-phi17*/	4, 33, 0, 2, 33, 1, 5, 98, 0, 1, 104, 1, 8, 
/* out0355_had-eta15-phi17*/	3, 33, 1, 5, 98, 0, 6, 98, 2, 2, 
/* out0356_had-eta16-phi17*/	2, 0, 0, 4, 98, 2, 7, 
/* out0357_had-eta17-phi17*/	4, 0, 0, 2, 0, 2, 3, 98, 2, 3, 102, 0, 2, 
/* out0358_had-eta18-phi17*/	3, 0, 2, 4, 102, 0, 1, 102, 1, 5, 
/* out0359_had-eta19-phi17*/	1, 102, 1, 5, 
/* out0360_had-eta0-phi18*/	1, 171, 0, 3, 
/* out0361_had-eta1-phi18*/	1, 171, 0, 4, 
/* out0362_had-eta2-phi18*/	2, 170, 0, 4, 171, 0, 1, 
/* out0363_had-eta3-phi18*/	1, 170, 0, 4, 
/* out0364_had-eta4-phi18*/	1, 169, 0, 4, 
/* out0365_had-eta5-phi18*/	5, 21, 0, 2, 23, 0, 6, 24, 0, 9, 24, 1, 16, 169, 0, 4, 
/* out0366_had-eta6-phi18*/	6, 20, 0, 4, 21, 2, 6, 23, 0, 3, 23, 1, 16, 23, 2, 1, 168, 0, 3, 
/* out0367_had-eta7-phi18*/	4, 20, 0, 8, 20, 1, 2, 20, 2, 13, 168, 0, 3, 
/* out0368_had-eta8-phi18*/	6, 16, 2, 1, 19, 0, 8, 19, 1, 5, 20, 1, 1, 20, 2, 3, 168, 0, 2, 
/* out0369_had-eta9-phi18*/	3, 15, 0, 5, 16, 2, 1, 19, 1, 11, 
/* out0370_had-eta10-phi18*/	2, 15, 0, 3, 15, 2, 10, 
/* out0371_had-eta11-phi18*/	4, 14, 0, 6, 15, 2, 5, 101, 0, 8, 101, 1, 3, 
/* out0372_had-eta12-phi18*/	5, 14, 0, 2, 14, 1, 7, 99, 0, 1, 101, 0, 1, 101, 1, 12, 
/* out0373_had-eta13-phi18*/	5, 1, 0, 2, 14, 1, 5, 99, 0, 6, 99, 2, 5, 101, 1, 1, 
/* out0374_had-eta14-phi18*/	4, 1, 0, 2, 1, 2, 5, 98, 0, 1, 99, 2, 8, 
/* out0375_had-eta15-phi18*/	4, 0, 0, 1, 1, 2, 5, 98, 0, 7, 98, 1, 2, 
/* out0376_had-eta16-phi18*/	2, 0, 0, 4, 98, 1, 6, 
/* out0377_had-eta17-phi18*/	4, 0, 0, 2, 0, 1, 2, 98, 1, 3, 128, 0, 2, 
/* out0378_had-eta18-phi18*/	3, 0, 1, 4, 128, 0, 1, 128, 2, 5, 
/* out0379_had-eta19-phi18*/	1, 128, 2, 5, 
/* out0380_had-eta0-phi19*/	1, 171, 0, 3, 
/* out0381_had-eta1-phi19*/	1, 171, 0, 4, 
/* out0382_had-eta2-phi19*/	2, 170, 0, 4, 171, 0, 1, 
/* out0383_had-eta3-phi19*/	1, 170, 0, 4, 
/* out0384_had-eta4-phi19*/	1, 169, 0, 4, 
/* out0385_had-eta5-phi19*/	6, 21, 0, 12, 21, 1, 1, 22, 0, 1, 22, 1, 16, 24, 0, 7, 169, 0, 4, 
/* out0386_had-eta6-phi19*/	6, 17, 0, 2, 20, 0, 1, 21, 0, 2, 21, 1, 12, 21, 2, 10, 168, 0, 3, 
/* out0387_had-eta7-phi19*/	6, 16, 0, 1, 17, 0, 1, 17, 2, 8, 20, 0, 3, 20, 1, 11, 168, 0, 3, 
/* out0388_had-eta8-phi19*/	5, 16, 0, 11, 16, 1, 1, 16, 2, 5, 20, 1, 2, 168, 0, 2, 
/* out0389_had-eta9-phi19*/	3, 15, 0, 5, 16, 1, 1, 16, 2, 9, 
/* out0390_had-eta10-phi19*/	2, 15, 0, 3, 15, 1, 10, 
/* out0391_had-eta11-phi19*/	6, 2, 0, 4, 2, 2, 1, 15, 1, 5, 15, 2, 1, 100, 0, 9, 100, 2, 4, 
/* out0392_had-eta12-phi19*/	4, 2, 2, 7, 14, 1, 3, 99, 0, 2, 100, 2, 11, 
/* out0393_had-eta13-phi19*/	5, 1, 0, 6, 2, 2, 1, 14, 1, 1, 99, 0, 7, 99, 1, 4, 
/* out0394_had-eta14-phi19*/	5, 1, 0, 4, 1, 1, 1, 1, 2, 1, 99, 1, 7, 99, 2, 2, 
/* out0395_had-eta15-phi19*/	7, 1, 1, 2, 1, 2, 4, 98, 0, 1, 98, 1, 2, 99, 2, 1, 129, 0, 2, 129, 2, 3, 
/* out0396_had-eta16-phi19*/	6, 0, 0, 2, 0, 1, 1, 1, 1, 1, 1, 2, 1, 98, 1, 3, 129, 2, 3, 
/* out0397_had-eta17-phi19*/	2, 0, 1, 5, 128, 0, 5, 
/* out0398_had-eta18-phi19*/	3, 0, 1, 4, 128, 0, 3, 128, 2, 2, 
/* out0399_had-eta19-phi19*/	1, 128, 2, 4, 
/* out0400_had-eta0-phi20*/	1, 175, 0, 3, 
/* out0401_had-eta1-phi20*/	1, 175, 0, 4, 
/* out0402_had-eta2-phi20*/	2, 174, 0, 4, 175, 0, 1, 
/* out0403_had-eta3-phi20*/	1, 174, 0, 4, 
/* out0404_had-eta4-phi20*/	2, 22, 0, 1, 173, 0, 4, 
/* out0405_had-eta5-phi20*/	6, 18, 0, 14, 18, 1, 1, 18, 2, 3, 21, 1, 1, 22, 0, 14, 173, 0, 4, 
/* out0406_had-eta6-phi20*/	6, 17, 0, 10, 17, 1, 1, 18, 1, 2, 18, 2, 13, 21, 1, 2, 172, 0, 3, 
/* out0407_had-eta7-phi20*/	5, 4, 0, 1, 17, 0, 3, 17, 1, 12, 17, 2, 7, 172, 0, 3, 
/* out0408_had-eta8-phi20*/	6, 4, 0, 2, 4, 2, 5, 16, 0, 4, 16, 1, 8, 17, 2, 1, 172, 0, 2, 
/* out0409_had-eta9-phi20*/	4, 3, 0, 9, 3, 2, 1, 4, 2, 1, 16, 1, 6, 
/* out0410_had-eta10-phi20*/	3, 3, 0, 1, 3, 2, 11, 15, 1, 1, 
/* out0411_had-eta11-phi20*/	6, 2, 0, 10, 2, 1, 1, 3, 2, 1, 100, 0, 7, 100, 1, 6, 131, 1, 1, 
/* out0412_had-eta12-phi20*/	6, 2, 0, 1, 2, 1, 4, 2, 2, 4, 100, 1, 10, 100, 2, 1, 130, 0, 3, 
/* out0413_had-eta13-phi20*/	7, 1, 0, 2, 1, 1, 1, 2, 1, 1, 2, 2, 3, 99, 1, 3, 130, 0, 2, 130, 2, 6, 
/* out0414_had-eta14-phi20*/	4, 1, 1, 6, 99, 1, 2, 129, 0, 5, 130, 2, 3, 
/* out0415_had-eta15-phi20*/	4, 1, 1, 5, 7, 0, 1, 129, 0, 5, 129, 2, 2, 
/* out0416_had-eta16-phi20*/	3, 7, 0, 3, 7, 2, 1, 129, 2, 6, 
/* out0417_had-eta17-phi20*/	4, 7, 2, 4, 128, 0, 4, 128, 1, 1, 129, 2, 1, 
/* out0418_had-eta18-phi20*/	3, 7, 2, 2, 128, 0, 1, 128, 1, 5, 
/* out0419_had-eta19-phi20*/	1, 128, 1, 3, 
/* out0420_had-eta0-phi21*/	1, 175, 0, 3, 
/* out0421_had-eta1-phi21*/	1, 175, 0, 4, 
/* out0422_had-eta2-phi21*/	2, 174, 0, 4, 175, 0, 1, 
/* out0423_had-eta3-phi21*/	1, 174, 0, 4, 
/* out0424_had-eta4-phi21*/	1, 173, 0, 4, 
/* out0425_had-eta5-phi21*/	5, 6, 0, 9, 6, 2, 9, 18, 0, 2, 18, 1, 6, 173, 0, 4, 
/* out0426_had-eta6-phi21*/	6, 5, 0, 14, 5, 1, 1, 5, 2, 4, 6, 2, 3, 18, 1, 7, 172, 0, 3, 
/* out0427_had-eta7-phi21*/	5, 4, 0, 8, 5, 1, 1, 5, 2, 12, 17, 1, 3, 172, 0, 3, 
/* out0428_had-eta8-phi21*/	4, 4, 0, 5, 4, 1, 7, 4, 2, 7, 172, 0, 2, 
/* out0429_had-eta9-phi21*/	5, 3, 0, 6, 3, 1, 4, 4, 1, 1, 4, 2, 3, 10, 2, 1, 
/* out0430_had-eta10-phi21*/	3, 3, 1, 10, 3, 2, 2, 9, 0, 1, 
/* out0431_had-eta11-phi21*/	8, 2, 0, 1, 2, 1, 3, 3, 1, 1, 3, 2, 1, 9, 0, 2, 9, 2, 3, 131, 0, 1, 131, 1, 9, 
/* out0432_had-eta12-phi21*/	5, 2, 1, 6, 8, 0, 2, 9, 2, 2, 130, 0, 8, 131, 1, 5, 
/* out0433_had-eta13-phi21*/	6, 2, 1, 1, 8, 0, 6, 8, 2, 1, 130, 0, 3, 130, 1, 5, 130, 2, 3, 
/* out0434_had-eta14-phi21*/	4, 8, 2, 6, 129, 0, 3, 130, 1, 2, 130, 2, 4, 
/* out0435_had-eta15-phi21*/	4, 7, 0, 4, 8, 2, 2, 129, 0, 1, 129, 1, 7, 
/* out0436_had-eta16-phi21*/	2, 7, 0, 4, 129, 1, 6, 
/* out0437_had-eta17-phi21*/	6, 7, 2, 4, 95, 0, 2, 95, 2, 2, 128, 1, 1, 129, 1, 1, 129, 2, 1, 
/* out0438_had-eta18-phi21*/	3, 7, 2, 3, 95, 2, 2, 128, 1, 4, 
/* out0439_had-eta19-phi21*/	1, 128, 1, 2, 
/* out0440_had-eta0-phi22*/	1, 179, 0, 3, 
/* out0441_had-eta1-phi22*/	1, 179, 0, 4, 
/* out0442_had-eta2-phi22*/	2, 178, 0, 4, 179, 0, 1, 
/* out0443_had-eta3-phi22*/	1, 178, 0, 4, 
/* out0444_had-eta4-phi22*/	1, 177, 0, 4, 
/* out0445_had-eta5-phi22*/	6, 6, 0, 7, 6, 1, 14, 6, 2, 2, 12, 0, 3, 13, 1, 7, 177, 0, 4, 
/* out0446_had-eta6-phi22*/	7, 5, 0, 2, 5, 1, 7, 6, 1, 2, 6, 2, 2, 12, 0, 5, 12, 2, 9, 176, 0, 3, 
/* out0447_had-eta7-phi22*/	5, 4, 1, 1, 5, 1, 7, 11, 0, 11, 11, 2, 4, 176, 0, 3, 
/* out0448_had-eta8-phi22*/	4, 4, 1, 7, 10, 0, 5, 11, 2, 8, 176, 0, 2, 
/* out0449_had-eta9-phi22*/	3, 10, 0, 8, 10, 1, 1, 10, 2, 8, 
/* out0450_had-eta10-phi22*/	3, 3, 1, 1, 9, 0, 7, 10, 2, 5, 
/* out0451_had-eta11-phi22*/	5, 9, 0, 5, 9, 1, 2, 9, 2, 4, 97, 0, 1, 131, 0, 10, 
/* out0452_had-eta12-phi22*/	7, 8, 0, 3, 9, 2, 6, 97, 0, 5, 97, 2, 4, 130, 1, 2, 131, 0, 5, 131, 1, 1, 
/* out0453_had-eta13-phi22*/	5, 8, 0, 5, 8, 1, 2, 96, 0, 2, 97, 2, 4, 130, 1, 6, 
/* out0454_had-eta14-phi22*/	5, 8, 1, 3, 8, 2, 4, 96, 0, 7, 96, 2, 2, 130, 1, 1, 
/* out0455_had-eta15-phi22*/	4, 7, 0, 2, 8, 2, 3, 96, 2, 7, 129, 1, 1, 
/* out0456_had-eta16-phi22*/	5, 7, 0, 2, 7, 1, 3, 95, 0, 5, 96, 2, 1, 129, 1, 1, 
/* out0457_had-eta17-phi22*/	3, 7, 1, 4, 95, 0, 4, 95, 2, 2, 
/* out0458_had-eta18-phi22*/	3, 7, 1, 2, 7, 2, 1, 95, 2, 5, 
/* out0459_had-eta19-phi22*/	2, 7, 2, 1, 95, 2, 1, 
/* out0460_had-eta0-phi23*/	1, 179, 0, 3, 
/* out0461_had-eta1-phi23*/	1, 179, 0, 4, 
/* out0462_had-eta2-phi23*/	2, 178, 0, 4, 179, 0, 1, 
/* out0463_had-eta3-phi23*/	1, 178, 0, 4, 
/* out0464_had-eta4-phi23*/	1, 177, 0, 4, 
/* out0465_had-eta5-phi23*/	5, 12, 0, 5, 12, 1, 1, 13, 0, 16, 13, 1, 9, 177, 0, 4, 
/* out0466_had-eta6-phi23*/	4, 12, 0, 3, 12, 1, 15, 12, 2, 6, 176, 0, 3, 
/* out0467_had-eta7-phi23*/	4, 11, 0, 5, 11, 1, 11, 12, 2, 1, 176, 0, 3, 
/* out0468_had-eta8-phi23*/	5, 10, 0, 2, 10, 1, 1, 11, 1, 5, 11, 2, 4, 176, 0, 2, 
/* out0469_had-eta9-phi23*/	2, 10, 0, 1, 10, 1, 12, 
/* out0470_had-eta10-phi23*/	4, 9, 0, 1, 9, 1, 2, 10, 1, 2, 10, 2, 2, 
/* out0471_had-eta11-phi23*/	3, 9, 1, 9, 97, 0, 5, 97, 1, 1, 
/* out0472_had-eta12-phi23*/	5, 9, 1, 3, 9, 2, 1, 97, 0, 5, 97, 1, 13, 97, 2, 2, 
/* out0473_had-eta13-phi23*/	5, 8, 1, 5, 96, 0, 3, 96, 1, 1, 97, 1, 2, 97, 2, 6, 
/* out0474_had-eta14-phi23*/	3, 8, 1, 5, 96, 0, 4, 96, 1, 5, 
/* out0475_had-eta15-phi23*/	3, 8, 1, 1, 96, 1, 4, 96, 2, 5, 
/* out0476_had-eta16-phi23*/	5, 7, 1, 3, 95, 0, 4, 95, 1, 7, 96, 1, 6, 96, 2, 1, 
/* out0477_had-eta17-phi23*/	3, 7, 1, 3, 95, 0, 1, 95, 1, 5, 
/* out0478_had-eta18-phi23*/	3, 7, 1, 1, 95, 1, 3, 95, 2, 2, 
/* out0479_had-eta19-phi23*/	2, 95, 1, 1, 95, 2, 2, 
};