parameter integer matrixH [0:4485] = {
/* num inputs = 156(in0-in155) */
/* num outputs = 560(out0-out559) */
//* max inputs per outputs = 8 */
//* total number of input in adders 1335 */

/* out0000_had-eta0-phi0*/	0, 
/* out0001_had-eta1-phi0*/	0, 
/* out0002_had-eta2-phi0*/	0, 
/* out0003_had-eta3-phi0*/	0, 
/* out0004_had-eta4-phi0*/	0, 
/* out0005_had-eta5-phi0*/	0, 
/* out0006_had-eta6-phi0*/	0, 
/* out0007_had-eta7-phi0*/	0, 
/* out0008_had-eta8-phi0*/	0, 
/* out0009_had-eta9-phi0*/	0, 
/* out0010_had-eta10-phi0*/	0, 
/* out0011_had-eta11-phi0*/	0, 
/* out0012_had-eta12-phi0*/	0, 
/* out0013_had-eta13-phi0*/	0, 
/* out0014_had-eta14-phi0*/	0, 
/* out0015_had-eta15-phi0*/	0, 
/* out0016_had-eta16-phi0*/	0, 
/* out0017_had-eta17-phi0*/	0, 
/* out0018_had-eta18-phi0*/	0, 
/* out0019_had-eta19-phi0*/	0, 
/* out0020_had-eta0-phi1*/	0, 
/* out0021_had-eta1-phi1*/	0, 
/* out0022_had-eta2-phi1*/	0, 
/* out0023_had-eta3-phi1*/	0, 
/* out0024_had-eta4-phi1*/	0, 
/* out0025_had-eta5-phi1*/	0, 
/* out0026_had-eta6-phi1*/	0, 
/* out0027_had-eta7-phi1*/	0, 
/* out0028_had-eta8-phi1*/	0, 
/* out0029_had-eta9-phi1*/	0, 
/* out0030_had-eta10-phi1*/	0, 
/* out0031_had-eta11-phi1*/	0, 
/* out0032_had-eta12-phi1*/	0, 
/* out0033_had-eta13-phi1*/	0, 
/* out0034_had-eta14-phi1*/	0, 
/* out0035_had-eta15-phi1*/	0, 
/* out0036_had-eta16-phi1*/	0, 
/* out0037_had-eta17-phi1*/	0, 
/* out0038_had-eta18-phi1*/	0, 
/* out0039_had-eta19-phi1*/	0, 
/* out0040_had-eta0-phi2*/	0, 
/* out0041_had-eta1-phi2*/	0, 
/* out0042_had-eta2-phi2*/	0, 
/* out0043_had-eta3-phi2*/	0, 
/* out0044_had-eta4-phi2*/	0, 
/* out0045_had-eta5-phi2*/	0, 
/* out0046_had-eta6-phi2*/	0, 
/* out0047_had-eta7-phi2*/	0, 
/* out0048_had-eta8-phi2*/	0, 
/* out0049_had-eta9-phi2*/	0, 
/* out0050_had-eta10-phi2*/	0, 
/* out0051_had-eta11-phi2*/	0, 
/* out0052_had-eta12-phi2*/	0, 
/* out0053_had-eta13-phi2*/	0, 
/* out0054_had-eta14-phi2*/	0, 
/* out0055_had-eta15-phi2*/	0, 
/* out0056_had-eta16-phi2*/	0, 
/* out0057_had-eta17-phi2*/	0, 
/* out0058_had-eta18-phi2*/	0, 
/* out0059_had-eta19-phi2*/	0, 
/* out0060_had-eta0-phi3*/	0, 
/* out0061_had-eta1-phi3*/	1, 133, 0, 1, 
/* out0062_had-eta2-phi3*/	2, 132, 0, 1, 133, 0, 7, 
/* out0063_had-eta3-phi3*/	1, 132, 0, 4, 
/* out0064_had-eta4-phi3*/	1, 132, 0, 3, 
/* out0065_had-eta5-phi3*/	3, 93, 2, 2, 94, 0, 4, 94, 1, 15, 
/* out0066_had-eta6-phi3*/	3, 93, 0, 1, 93, 1, 10, 93, 2, 13, 
/* out0067_had-eta7-phi3*/	2, 92, 2, 13, 93, 1, 4, 
/* out0068_had-eta8-phi3*/	2, 91, 2, 2, 92, 1, 12, 
/* out0069_had-eta9-phi3*/	2, 91, 1, 4, 91, 2, 9, 
/* out0070_had-eta10-phi3*/	2, 90, 2, 2, 91, 1, 6, 
/* out0071_had-eta11-phi3*/	3, 90, 1, 3, 90, 2, 7, 127, 1, 8, 
/* out0072_had-eta12-phi3*/	3, 90, 1, 5, 126, 2, 5, 127, 1, 2, 
/* out0073_had-eta13-phi3*/	3, 89, 2, 4, 126, 1, 5, 126, 2, 4, 
/* out0074_had-eta14-phi3*/	4, 89, 1, 4, 89, 2, 2, 125, 2, 1, 126, 1, 2, 
/* out0075_had-eta15-phi3*/	3, 89, 1, 1, 125, 1, 1, 125, 2, 5, 
/* out0076_had-eta16-phi3*/	2, 88, 2, 2, 125, 1, 4, 
/* out0077_had-eta17-phi3*/	3, 88, 1, 2, 88, 2, 2, 124, 1, 1, 
/* out0078_had-eta18-phi3*/	2, 88, 1, 1, 124, 1, 3, 
/* out0079_had-eta19-phi3*/	0, 
/* out0080_had-eta0-phi4*/	0, 
/* out0081_had-eta1-phi4*/	1, 133, 0, 1, 
/* out0082_had-eta2-phi4*/	2, 132, 0, 1, 133, 0, 7, 
/* out0083_had-eta3-phi4*/	1, 132, 0, 4, 
/* out0084_had-eta4-phi4*/	1, 132, 0, 3, 
/* out0085_had-eta5-phi4*/	5, 87, 1, 5, 87, 2, 15, 93, 2, 1, 94, 0, 12, 94, 1, 1, 
/* out0086_had-eta6-phi4*/	4, 86, 2, 7, 87, 1, 7, 93, 0, 14, 93, 1, 1, 
/* out0087_had-eta7-phi4*/	6, 86, 1, 7, 86, 2, 2, 92, 0, 9, 92, 2, 3, 93, 0, 1, 93, 1, 1, 
/* out0088_had-eta8-phi4*/	6, 85, 1, 2, 85, 2, 5, 91, 0, 1, 91, 2, 2, 92, 0, 7, 92, 1, 4, 
/* out0089_had-eta9-phi4*/	4, 85, 1, 1, 91, 0, 11, 91, 1, 1, 91, 2, 3, 
/* out0090_had-eta10-phi4*/	5, 84, 2, 1, 90, 0, 2, 90, 2, 3, 91, 0, 3, 91, 1, 5, 
/* out0091_had-eta11-phi4*/	6, 90, 0, 6, 90, 1, 1, 90, 2, 4, 122, 2, 1, 127, 0, 14, 127, 1, 4, 
/* out0092_had-eta12-phi4*/	8, 89, 2, 2, 90, 0, 1, 90, 1, 7, 122, 1, 1, 126, 0, 4, 126, 2, 6, 127, 0, 1, 127, 1, 2, 
/* out0093_had-eta13-phi4*/	5, 89, 0, 1, 89, 2, 7, 126, 0, 5, 126, 1, 5, 126, 2, 1, 
/* out0094_had-eta14-phi4*/	5, 89, 0, 1, 89, 1, 5, 89, 2, 1, 125, 2, 5, 126, 1, 4, 
/* out0095_had-eta15-phi4*/	5, 88, 2, 2, 89, 1, 4, 125, 0, 2, 125, 1, 1, 125, 2, 5, 
/* out0096_had-eta16-phi4*/	2, 88, 2, 5, 125, 1, 6, 
/* out0097_had-eta17-phi4*/	4, 88, 1, 2, 88, 2, 1, 124, 1, 4, 125, 1, 1, 
/* out0098_had-eta18-phi4*/	2, 88, 1, 3, 124, 1, 4, 
/* out0099_had-eta19-phi4*/	1, 88, 1, 1, 
/* out0100_had-eta0-phi5*/	0, 
/* out0101_had-eta1-phi5*/	1, 135, 0, 1, 
/* out0102_had-eta2-phi5*/	2, 134, 0, 1, 135, 0, 7, 
/* out0103_had-eta3-phi5*/	1, 134, 0, 4, 
/* out0104_had-eta4-phi5*/	1, 134, 0, 3, 
/* out0105_had-eta5-phi5*/	3, 81, 2, 5, 87, 0, 14, 87, 2, 1, 
/* out0106_had-eta6-phi5*/	6, 81, 1, 6, 81, 2, 4, 86, 0, 8, 86, 2, 6, 87, 0, 2, 87, 1, 4, 
/* out0107_had-eta7-phi5*/	7, 80, 1, 1, 80, 2, 2, 85, 0, 1, 85, 2, 3, 86, 0, 8, 86, 1, 9, 86, 2, 1, 
/* out0108_had-eta8-phi5*/	3, 85, 0, 7, 85, 1, 5, 85, 2, 8, 
/* out0109_had-eta9-phi5*/	3, 84, 2, 8, 85, 1, 7, 91, 0, 1, 
/* out0110_had-eta10-phi5*/	2, 84, 1, 8, 84, 2, 6, 
/* out0111_had-eta11-phi5*/	5, 83, 2, 3, 84, 1, 3, 90, 0, 5, 122, 2, 13, 127, 0, 1, 
/* out0112_had-eta12-phi5*/	6, 83, 1, 2, 83, 2, 4, 90, 0, 2, 122, 1, 10, 122, 2, 1, 126, 0, 2, 
/* out0113_had-eta13-phi5*/	4, 83, 1, 2, 89, 0, 7, 121, 2, 6, 126, 0, 5, 
/* out0114_had-eta14-phi5*/	4, 89, 0, 6, 121, 1, 4, 121, 2, 2, 125, 0, 2, 
/* out0115_had-eta15-phi5*/	6, 82, 2, 1, 88, 0, 1, 88, 2, 2, 89, 0, 1, 89, 1, 2, 125, 0, 7, 
/* out0116_had-eta16-phi5*/	5, 88, 0, 3, 88, 2, 2, 120, 2, 1, 125, 0, 4, 125, 1, 2, 
/* out0117_had-eta17-phi5*/	5, 88, 0, 2, 88, 1, 2, 124, 0, 3, 124, 1, 3, 125, 1, 1, 
/* out0118_had-eta18-phi5*/	3, 88, 1, 3, 124, 0, 5, 124, 1, 1, 
/* out0119_had-eta19-phi5*/	1, 88, 1, 1, 
/* out0120_had-eta0-phi6*/	0, 
/* out0121_had-eta1-phi6*/	1, 135, 0, 1, 
/* out0122_had-eta2-phi6*/	2, 134, 0, 1, 135, 0, 7, 
/* out0123_had-eta3-phi6*/	1, 134, 0, 4, 
/* out0124_had-eta4-phi6*/	1, 134, 0, 3, 
/* out0125_had-eta5-phi6*/	4, 76, 1, 7, 76, 2, 16, 81, 0, 8, 81, 2, 6, 
/* out0126_had-eta6-phi6*/	7, 75, 1, 1, 75, 2, 2, 80, 0, 2, 80, 2, 5, 81, 0, 8, 81, 1, 10, 81, 2, 1, 
/* out0127_had-eta7-phi6*/	3, 80, 0, 5, 80, 1, 9, 80, 2, 9, 
/* out0128_had-eta8-phi6*/	3, 79, 2, 9, 80, 1, 4, 85, 0, 7, 
/* out0129_had-eta9-phi6*/	6, 79, 1, 6, 79, 2, 2, 84, 0, 6, 84, 2, 1, 85, 0, 1, 85, 1, 1, 
/* out0130_had-eta10-phi6*/	3, 78, 2, 1, 84, 0, 10, 84, 1, 3, 
/* out0131_had-eta11-phi6*/	5, 83, 0, 3, 83, 2, 6, 84, 1, 2, 122, 0, 11, 122, 2, 1, 
/* out0132_had-eta12-phi6*/	7, 83, 0, 2, 83, 1, 4, 83, 2, 3, 121, 2, 1, 122, 0, 5, 122, 1, 5, 123, 2, 1, 
/* out0133_had-eta13-phi6*/	4, 82, 2, 2, 83, 1, 6, 121, 0, 4, 121, 2, 7, 
/* out0134_had-eta14-phi6*/	3, 82, 2, 6, 121, 0, 1, 121, 1, 8, 
/* out0135_had-eta15-phi6*/	5, 82, 1, 4, 82, 2, 1, 120, 2, 4, 121, 1, 2, 125, 0, 1, 
/* out0136_had-eta16-phi6*/	4, 82, 1, 1, 88, 0, 4, 120, 1, 1, 120, 2, 5, 
/* out0137_had-eta17-phi6*/	3, 88, 0, 4, 120, 1, 4, 124, 0, 3, 
/* out0138_had-eta18-phi6*/	3, 88, 0, 2, 88, 1, 1, 124, 0, 5, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	0, 
/* out0141_had-eta1-phi7*/	1, 137, 0, 1, 
/* out0142_had-eta2-phi7*/	2, 136, 0, 1, 137, 0, 7, 
/* out0143_had-eta3-phi7*/	1, 136, 0, 4, 
/* out0144_had-eta4-phi7*/	1, 136, 0, 3, 
/* out0145_had-eta5-phi7*/	6, 75, 0, 3, 75, 2, 5, 76, 0, 16, 76, 1, 9, 77, 1, 2, 77, 2, 11, 
/* out0146_had-eta6-phi7*/	3, 75, 0, 6, 75, 1, 13, 75, 2, 9, 
/* out0147_had-eta7-phi7*/	5, 74, 1, 2, 74, 2, 11, 75, 1, 1, 80, 0, 9, 80, 1, 1, 
/* out0148_had-eta8-phi7*/	4, 74, 1, 4, 79, 0, 11, 79, 2, 5, 80, 1, 1, 
/* out0149_had-eta9-phi7*/	3, 78, 2, 3, 79, 0, 4, 79, 1, 10, 
/* out0150_had-eta10-phi7*/	2, 78, 1, 2, 78, 2, 12, 
/* out0151_had-eta11-phi7*/	3, 78, 1, 7, 83, 0, 4, 123, 2, 9, 
/* out0152_had-eta12-phi7*/	4, 63, 2, 2, 83, 0, 7, 123, 1, 7, 123, 2, 6, 
/* out0153_had-eta13-phi7*/	7, 63, 2, 1, 82, 0, 2, 82, 2, 3, 83, 1, 2, 116, 2, 1, 121, 0, 7, 123, 1, 3, 
/* out0154_had-eta14-phi7*/	5, 82, 0, 3, 82, 2, 3, 116, 2, 2, 121, 0, 4, 121, 1, 2, 
/* out0155_had-eta15-phi7*/	3, 82, 1, 5, 120, 0, 3, 120, 2, 4, 
/* out0156_had-eta16-phi7*/	5, 49, 2, 2, 82, 1, 3, 120, 0, 2, 120, 1, 2, 120, 2, 2, 
/* out0157_had-eta17-phi7*/	2, 49, 2, 3, 120, 1, 5, 
/* out0158_had-eta18-phi7*/	3, 49, 1, 2, 49, 2, 2, 120, 1, 1, 
/* out0159_had-eta19-phi7*/	0, 
/* out0160_had-eta0-phi8*/	0, 
/* out0161_had-eta1-phi8*/	1, 137, 0, 1, 
/* out0162_had-eta2-phi8*/	2, 136, 0, 1, 137, 0, 7, 
/* out0163_had-eta3-phi8*/	1, 136, 0, 4, 
/* out0164_had-eta4-phi8*/	1, 136, 0, 3, 
/* out0165_had-eta5-phi8*/	5, 70, 2, 3, 75, 0, 1, 77, 0, 16, 77, 1, 14, 77, 2, 5, 
/* out0166_had-eta6-phi8*/	6, 70, 1, 6, 70, 2, 13, 74, 0, 1, 74, 2, 1, 75, 0, 6, 75, 1, 1, 
/* out0167_had-eta7-phi8*/	4, 70, 1, 1, 74, 0, 15, 74, 1, 3, 74, 2, 4, 
/* out0168_had-eta8-phi8*/	3, 68, 2, 10, 74, 1, 7, 79, 0, 1, 
/* out0169_had-eta9-phi8*/	3, 68, 1, 7, 68, 2, 6, 78, 0, 2, 
/* out0170_had-eta10-phi8*/	2, 78, 0, 13, 78, 1, 1, 
/* out0171_had-eta11-phi8*/	4, 63, 2, 4, 78, 0, 1, 78, 1, 6, 123, 0, 8, 
/* out0172_had-eta12-phi8*/	4, 63, 1, 1, 63, 2, 9, 123, 0, 8, 123, 1, 4, 
/* out0173_had-eta13-phi8*/	4, 63, 1, 6, 82, 0, 1, 116, 2, 8, 123, 1, 2, 
/* out0174_had-eta14-phi8*/	3, 82, 0, 7, 116, 1, 4, 116, 2, 5, 
/* out0175_had-eta15-phi8*/	4, 82, 0, 3, 82, 1, 2, 116, 1, 3, 120, 0, 4, 
/* out0176_had-eta16-phi8*/	3, 49, 2, 4, 82, 1, 1, 120, 0, 6, 
/* out0177_had-eta17-phi8*/	3, 49, 2, 4, 120, 0, 1, 120, 1, 3, 
/* out0178_had-eta18-phi8*/	2, 49, 1, 5, 49, 2, 1, 
/* out0179_had-eta19-phi8*/	1, 49, 1, 1, 
/* out0180_had-eta0-phi9*/	0, 
/* out0181_had-eta1-phi9*/	1, 139, 0, 1, 
/* out0182_had-eta2-phi9*/	2, 138, 0, 1, 139, 0, 7, 
/* out0183_had-eta3-phi9*/	1, 138, 0, 4, 
/* out0184_had-eta4-phi9*/	1, 138, 0, 3, 
/* out0185_had-eta5-phi9*/	5, 70, 0, 3, 71, 2, 1, 72, 0, 5, 72, 1, 14, 72, 2, 16, 
/* out0186_had-eta6-phi9*/	6, 69, 0, 1, 69, 2, 1, 70, 0, 13, 70, 1, 7, 71, 1, 1, 71, 2, 6, 
/* out0187_had-eta7-phi9*/	4, 69, 0, 4, 69, 1, 3, 69, 2, 15, 70, 1, 2, 
/* out0188_had-eta8-phi9*/	3, 65, 2, 1, 68, 0, 11, 69, 1, 7, 
/* out0189_had-eta9-phi9*/	3, 64, 2, 2, 68, 0, 5, 68, 1, 8, 
/* out0190_had-eta10-phi9*/	3, 64, 1, 1, 64, 2, 13, 68, 1, 1, 
/* out0191_had-eta11-phi9*/	4, 63, 0, 5, 64, 1, 6, 64, 2, 1, 118, 2, 8, 
/* out0192_had-eta12-phi9*/	4, 63, 0, 8, 63, 1, 1, 118, 1, 4, 118, 2, 8, 
/* out0193_had-eta13-phi9*/	4, 50, 2, 1, 63, 1, 7, 116, 0, 8, 118, 1, 2, 
/* out0194_had-eta14-phi9*/	3, 50, 2, 7, 116, 0, 5, 116, 1, 4, 
/* out0195_had-eta15-phi9*/	4, 50, 1, 2, 50, 2, 3, 115, 2, 4, 116, 1, 4, 
/* out0196_had-eta16-phi9*/	3, 49, 0, 4, 50, 1, 1, 115, 2, 6, 
/* out0197_had-eta17-phi9*/	3, 49, 0, 4, 115, 1, 3, 115, 2, 1, 
/* out0198_had-eta18-phi9*/	1, 49, 1, 5, 
/* out0199_had-eta19-phi9*/	1, 49, 1, 1, 
/* out0200_had-eta0-phi10*/	0, 
/* out0201_had-eta1-phi10*/	1, 139, 0, 1, 
/* out0202_had-eta2-phi10*/	2, 138, 0, 1, 139, 0, 7, 
/* out0203_had-eta3-phi10*/	1, 138, 0, 4, 
/* out0204_had-eta4-phi10*/	1, 138, 0, 3, 
/* out0205_had-eta5-phi10*/	6, 71, 0, 5, 71, 2, 3, 72, 0, 11, 72, 1, 2, 73, 1, 9, 73, 2, 16, 
/* out0206_had-eta6-phi10*/	3, 71, 0, 9, 71, 1, 13, 71, 2, 6, 
/* out0207_had-eta7-phi10*/	5, 66, 1, 1, 66, 2, 9, 69, 0, 11, 69, 1, 2, 71, 1, 1, 
/* out0208_had-eta8-phi10*/	4, 65, 0, 5, 65, 2, 11, 66, 1, 1, 69, 1, 4, 
/* out0209_had-eta9-phi10*/	3, 64, 0, 3, 65, 1, 10, 65, 2, 4, 
/* out0210_had-eta10-phi10*/	2, 64, 0, 12, 64, 1, 2, 
/* out0211_had-eta11-phi10*/	3, 51, 2, 4, 64, 1, 7, 118, 0, 9, 
/* out0212_had-eta12-phi10*/	4, 51, 2, 7, 63, 0, 2, 118, 0, 6, 118, 1, 7, 
/* out0213_had-eta13-phi10*/	8, 50, 0, 3, 50, 2, 2, 51, 1, 2, 63, 0, 1, 63, 1, 1, 116, 0, 1, 117, 2, 7, 118, 1, 3, 
/* out0214_had-eta14-phi10*/	6, 50, 0, 3, 50, 2, 3, 116, 0, 2, 116, 1, 1, 117, 1, 2, 117, 2, 4, 
/* out0215_had-eta15-phi10*/	3, 50, 1, 5, 115, 0, 4, 115, 2, 3, 
/* out0216_had-eta16-phi10*/	5, 49, 0, 2, 50, 1, 3, 115, 0, 2, 115, 1, 2, 115, 2, 2, 
/* out0217_had-eta17-phi10*/	2, 49, 0, 4, 115, 1, 5, 
/* out0218_had-eta18-phi10*/	3, 49, 0, 2, 49, 1, 2, 115, 1, 1, 
/* out0219_had-eta19-phi10*/	0, 
/* out0220_had-eta0-phi11*/	0, 
/* out0221_had-eta1-phi11*/	1, 141, 0, 1, 
/* out0222_had-eta2-phi11*/	2, 140, 0, 1, 141, 0, 7, 
/* out0223_had-eta3-phi11*/	1, 140, 0, 4, 
/* out0224_had-eta4-phi11*/	1, 140, 0, 3, 
/* out0225_had-eta5-phi11*/	4, 67, 0, 6, 67, 2, 8, 73, 0, 16, 73, 1, 7, 
/* out0226_had-eta6-phi11*/	7, 66, 0, 5, 66, 2, 2, 67, 0, 1, 67, 1, 10, 67, 2, 8, 71, 0, 2, 71, 1, 1, 
/* out0227_had-eta7-phi11*/	3, 66, 0, 9, 66, 1, 9, 66, 2, 5, 
/* out0228_had-eta8-phi11*/	3, 53, 2, 7, 65, 0, 9, 66, 1, 4, 
/* out0229_had-eta9-phi11*/	6, 52, 0, 1, 52, 2, 6, 53, 1, 1, 53, 2, 1, 65, 0, 2, 65, 1, 6, 
/* out0230_had-eta10-phi11*/	3, 52, 1, 3, 52, 2, 10, 64, 0, 1, 
/* out0231_had-eta11-phi11*/	5, 51, 0, 6, 51, 2, 3, 52, 1, 2, 119, 0, 1, 119, 2, 11, 
/* out0232_had-eta12-phi11*/	7, 51, 0, 3, 51, 1, 4, 51, 2, 2, 117, 0, 1, 118, 0, 1, 119, 1, 5, 119, 2, 5, 
/* out0233_had-eta13-phi11*/	4, 50, 0, 2, 51, 1, 6, 117, 0, 7, 117, 2, 4, 
/* out0234_had-eta14-phi11*/	3, 50, 0, 6, 117, 1, 8, 117, 2, 1, 
/* out0235_had-eta15-phi11*/	5, 50, 0, 1, 50, 1, 4, 112, 2, 1, 115, 0, 4, 117, 1, 2, 
/* out0236_had-eta16-phi11*/	4, 50, 1, 1, 56, 2, 4, 115, 0, 5, 115, 1, 1, 
/* out0237_had-eta17-phi11*/	3, 56, 2, 4, 111, 1, 3, 115, 1, 4, 
/* out0238_had-eta18-phi11*/	3, 56, 1, 1, 56, 2, 2, 111, 1, 5, 
/* out0239_had-eta19-phi11*/	0, 
/* out0240_had-eta0-phi12*/	0, 
/* out0241_had-eta1-phi12*/	1, 141, 0, 1, 
/* out0242_had-eta2-phi12*/	2, 140, 0, 1, 141, 0, 7, 
/* out0243_had-eta3-phi12*/	1, 140, 0, 4, 
/* out0244_had-eta4-phi12*/	1, 140, 0, 3, 
/* out0245_had-eta5-phi12*/	3, 55, 0, 1, 55, 2, 14, 67, 0, 5, 
/* out0246_had-eta6-phi12*/	6, 54, 0, 6, 54, 2, 8, 55, 1, 4, 55, 2, 2, 67, 0, 4, 67, 1, 6, 
/* out0247_had-eta7-phi12*/	7, 53, 0, 3, 53, 2, 1, 54, 0, 1, 54, 1, 9, 54, 2, 8, 66, 0, 2, 66, 1, 1, 
/* out0248_had-eta8-phi12*/	3, 53, 0, 8, 53, 1, 5, 53, 2, 7, 
/* out0249_had-eta9-phi12*/	3, 52, 0, 8, 53, 1, 7, 59, 2, 1, 
/* out0250_had-eta10-phi12*/	2, 52, 0, 6, 52, 1, 8, 
/* out0251_had-eta11-phi12*/	5, 51, 0, 3, 52, 1, 3, 58, 2, 5, 114, 1, 1, 119, 0, 13, 
/* out0252_had-eta12-phi12*/	6, 51, 0, 4, 51, 1, 2, 58, 2, 2, 113, 2, 2, 119, 0, 1, 119, 1, 10, 
/* out0253_had-eta13-phi12*/	4, 51, 1, 2, 57, 2, 7, 113, 2, 5, 117, 0, 6, 
/* out0254_had-eta14-phi12*/	4, 57, 2, 6, 112, 2, 2, 117, 0, 2, 117, 1, 4, 
/* out0255_had-eta15-phi12*/	6, 50, 0, 1, 56, 0, 2, 56, 2, 1, 57, 1, 2, 57, 2, 1, 112, 2, 7, 
/* out0256_had-eta16-phi12*/	5, 56, 0, 2, 56, 2, 3, 112, 1, 2, 112, 2, 4, 115, 0, 1, 
/* out0257_had-eta17-phi12*/	5, 56, 1, 2, 56, 2, 2, 111, 0, 3, 111, 1, 3, 112, 1, 1, 
/* out0258_had-eta18-phi12*/	3, 56, 1, 3, 111, 0, 1, 111, 1, 5, 
/* out0259_had-eta19-phi12*/	1, 56, 1, 1, 
/* out0260_had-eta0-phi13*/	0, 
/* out0261_had-eta1-phi13*/	1, 143, 0, 1, 
/* out0262_had-eta2-phi13*/	2, 142, 0, 1, 143, 0, 7, 
/* out0263_had-eta3-phi13*/	1, 142, 0, 4, 
/* out0264_had-eta4-phi13*/	1, 142, 0, 3, 
/* out0265_had-eta5-phi13*/	5, 55, 0, 15, 55, 1, 5, 61, 0, 1, 62, 0, 1, 62, 1, 12, 
/* out0266_had-eta6-phi13*/	4, 54, 0, 7, 55, 1, 7, 61, 1, 1, 61, 2, 14, 
/* out0267_had-eta7-phi13*/	6, 54, 0, 2, 54, 1, 7, 60, 0, 3, 60, 2, 9, 61, 1, 1, 61, 2, 1, 
/* out0268_had-eta8-phi13*/	6, 53, 0, 5, 53, 1, 2, 59, 0, 2, 59, 2, 1, 60, 1, 4, 60, 2, 7, 
/* out0269_had-eta9-phi13*/	4, 53, 1, 1, 59, 0, 3, 59, 1, 1, 59, 2, 11, 
/* out0270_had-eta10-phi13*/	5, 52, 0, 1, 58, 0, 4, 58, 2, 2, 59, 1, 5, 59, 2, 3, 
/* out0271_had-eta11-phi13*/	6, 58, 0, 4, 58, 1, 1, 58, 2, 6, 114, 0, 4, 114, 1, 14, 119, 0, 1, 
/* out0272_had-eta12-phi13*/	8, 57, 0, 2, 58, 1, 7, 58, 2, 1, 113, 0, 6, 113, 2, 4, 114, 0, 2, 114, 1, 1, 119, 1, 1, 
/* out0273_had-eta13-phi13*/	5, 57, 0, 7, 57, 2, 1, 113, 0, 1, 113, 1, 5, 113, 2, 5, 
/* out0274_had-eta14-phi13*/	5, 57, 0, 1, 57, 1, 5, 57, 2, 1, 112, 0, 5, 113, 1, 4, 
/* out0275_had-eta15-phi13*/	5, 56, 0, 2, 57, 1, 4, 112, 0, 5, 112, 1, 1, 112, 2, 2, 
/* out0276_had-eta16-phi13*/	2, 56, 0, 5, 112, 1, 6, 
/* out0277_had-eta17-phi13*/	4, 56, 0, 1, 56, 1, 2, 111, 0, 4, 112, 1, 1, 
/* out0278_had-eta18-phi13*/	2, 56, 1, 3, 111, 0, 4, 
/* out0279_had-eta19-phi13*/	1, 56, 1, 1, 
/* out0280_had-eta0-phi14*/	0, 
/* out0281_had-eta1-phi14*/	1, 143, 0, 1, 
/* out0282_had-eta2-phi14*/	2, 142, 0, 1, 143, 0, 7, 
/* out0283_had-eta3-phi14*/	1, 142, 0, 4, 
/* out0284_had-eta4-phi14*/	1, 142, 0, 3, 
/* out0285_had-eta5-phi14*/	4, 48, 2, 5, 61, 0, 2, 62, 0, 15, 62, 1, 4, 
/* out0286_had-eta6-phi14*/	5, 47, 2, 1, 48, 2, 3, 61, 0, 13, 61, 1, 10, 61, 2, 1, 
/* out0287_had-eta7-phi14*/	3, 47, 2, 6, 60, 0, 13, 61, 1, 4, 
/* out0288_had-eta8-phi14*/	3, 46, 2, 5, 59, 0, 2, 60, 1, 12, 
/* out0289_had-eta9-phi14*/	3, 46, 2, 2, 59, 0, 9, 59, 1, 4, 
/* out0290_had-eta10-phi14*/	3, 45, 2, 6, 58, 0, 2, 59, 1, 6, 
/* out0291_had-eta11-phi14*/	5, 45, 2, 2, 58, 0, 6, 58, 1, 3, 110, 2, 2, 114, 0, 8, 
/* out0292_had-eta12-phi14*/	5, 44, 2, 4, 58, 1, 5, 110, 2, 5, 113, 0, 5, 114, 0, 2, 
/* out0293_had-eta13-phi14*/	5, 44, 2, 3, 57, 0, 4, 109, 2, 1, 113, 0, 4, 113, 1, 5, 
/* out0294_had-eta14-phi14*/	6, 43, 2, 1, 57, 0, 2, 57, 1, 4, 109, 2, 5, 112, 0, 1, 113, 1, 2, 
/* out0295_had-eta15-phi14*/	5, 43, 2, 4, 57, 1, 1, 109, 2, 2, 112, 0, 5, 112, 1, 1, 
/* out0296_had-eta16-phi14*/	4, 43, 2, 3, 56, 0, 2, 108, 2, 2, 112, 1, 4, 
/* out0297_had-eta17-phi14*/	5, 42, 1, 1, 56, 0, 2, 56, 1, 2, 108, 2, 4, 111, 0, 1, 
/* out0298_had-eta18-phi14*/	4, 42, 1, 4, 56, 1, 1, 108, 2, 1, 111, 0, 3, 
/* out0299_had-eta19-phi14*/	1, 42, 1, 3, 
/* out0300_had-eta0-phi15*/	0, 
/* out0301_had-eta1-phi15*/	1, 145, 0, 1, 
/* out0302_had-eta2-phi15*/	2, 144, 0, 1, 145, 0, 7, 
/* out0303_had-eta3-phi15*/	1, 144, 0, 4, 
/* out0304_had-eta4-phi15*/	1, 144, 0, 3, 
/* out0305_had-eta5-phi15*/	4, 41, 1, 4, 48, 0, 15, 48, 1, 2, 48, 2, 5, 
/* out0306_had-eta6-phi15*/	5, 40, 2, 1, 47, 0, 10, 47, 2, 2, 48, 1, 13, 48, 2, 3, 
/* out0307_had-eta7-phi15*/	3, 47, 0, 4, 47, 1, 13, 47, 2, 7, 
/* out0308_had-eta8-phi15*/	3, 46, 0, 12, 46, 1, 2, 46, 2, 6, 
/* out0309_had-eta9-phi15*/	3, 45, 0, 4, 46, 1, 9, 46, 2, 3, 
/* out0310_had-eta10-phi15*/	3, 45, 0, 6, 45, 1, 2, 45, 2, 6, 
/* out0311_had-eta11-phi15*/	5, 44, 0, 3, 45, 1, 7, 45, 2, 2, 110, 0, 8, 110, 2, 2, 
/* out0312_had-eta12-phi15*/	5, 44, 0, 5, 44, 2, 5, 110, 0, 2, 110, 1, 5, 110, 2, 6, 
/* out0313_had-eta13-phi15*/	6, 44, 1, 4, 44, 2, 4, 109, 0, 5, 109, 2, 1, 110, 1, 4, 110, 2, 1, 
/* out0314_had-eta14-phi15*/	6, 43, 0, 4, 43, 2, 1, 44, 1, 2, 109, 0, 2, 109, 1, 1, 109, 2, 5, 
/* out0315_had-eta15-phi15*/	5, 43, 0, 1, 43, 2, 4, 108, 0, 1, 109, 1, 5, 109, 2, 2, 
/* out0316_had-eta16-phi15*/	4, 43, 1, 2, 43, 2, 3, 108, 0, 4, 108, 2, 3, 
/* out0317_had-eta17-phi15*/	5, 42, 0, 2, 42, 1, 1, 43, 1, 2, 108, 1, 1, 108, 2, 4, 
/* out0318_had-eta18-phi15*/	4, 42, 0, 1, 42, 1, 4, 108, 1, 3, 108, 2, 2, 
/* out0319_had-eta19-phi15*/	1, 42, 1, 3, 
/* out0320_had-eta0-phi16*/	0, 
/* out0321_had-eta1-phi16*/	1, 145, 0, 1, 
/* out0322_had-eta2-phi16*/	2, 144, 0, 1, 145, 0, 7, 
/* out0323_had-eta3-phi16*/	1, 144, 0, 4, 
/* out0324_had-eta4-phi16*/	1, 144, 0, 3, 
/* out0325_had-eta5-phi16*/	5, 40, 0, 5, 41, 0, 15, 41, 1, 12, 48, 0, 1, 48, 1, 1, 
/* out0326_had-eta6-phi16*/	4, 40, 0, 7, 40, 1, 7, 40, 2, 14, 47, 0, 1, 
/* out0327_had-eta7-phi16*/	6, 39, 0, 7, 39, 2, 9, 40, 1, 2, 40, 2, 1, 47, 0, 1, 47, 1, 3, 
/* out0328_had-eta8-phi16*/	6, 38, 0, 2, 38, 2, 1, 39, 1, 5, 39, 2, 7, 46, 0, 4, 46, 1, 2, 
/* out0329_had-eta9-phi16*/	4, 38, 0, 1, 38, 2, 11, 45, 0, 1, 46, 1, 3, 
/* out0330_had-eta10-phi16*/	5, 37, 2, 2, 38, 1, 1, 38, 2, 3, 45, 0, 5, 45, 1, 3, 
/* out0331_had-eta11-phi16*/	6, 37, 2, 6, 44, 0, 1, 45, 1, 4, 107, 0, 1, 107, 1, 14, 110, 0, 4, 
/* out0332_had-eta12-phi16*/	8, 37, 2, 1, 44, 0, 7, 44, 1, 2, 105, 0, 1, 105, 2, 4, 107, 1, 1, 110, 0, 2, 110, 1, 6, 
/* out0333_had-eta13-phi16*/	5, 36, 2, 1, 44, 1, 7, 105, 2, 5, 109, 0, 5, 110, 1, 1, 
/* out0334_had-eta14-phi16*/	5, 36, 2, 1, 43, 0, 5, 44, 1, 1, 109, 0, 4, 109, 1, 5, 
/* out0335_had-eta15-phi16*/	5, 43, 0, 4, 43, 1, 2, 103, 2, 2, 108, 0, 1, 109, 1, 5, 
/* out0336_had-eta16-phi16*/	2, 43, 1, 5, 108, 0, 6, 
/* out0337_had-eta17-phi16*/	4, 42, 0, 2, 43, 1, 1, 108, 0, 1, 108, 1, 4, 
/* out0338_had-eta18-phi16*/	2, 42, 0, 3, 108, 1, 4, 
/* out0339_had-eta19-phi16*/	1, 42, 0, 1, 
/* out0340_had-eta0-phi17*/	0, 
/* out0341_had-eta1-phi17*/	1, 147, 0, 1, 
/* out0342_had-eta2-phi17*/	2, 146, 0, 1, 147, 0, 7, 
/* out0343_had-eta3-phi17*/	1, 146, 0, 4, 
/* out0344_had-eta4-phi17*/	1, 146, 0, 3, 
/* out0345_had-eta5-phi17*/	4, 24, 0, 13, 24, 1, 5, 24, 2, 14, 41, 0, 1, 
/* out0346_had-eta6-phi17*/	6, 23, 0, 6, 23, 2, 8, 24, 1, 4, 24, 2, 2, 40, 0, 4, 40, 1, 6, 
/* out0347_had-eta7-phi17*/	7, 22, 0, 1, 22, 2, 1, 23, 1, 2, 23, 2, 8, 39, 0, 9, 39, 1, 3, 40, 1, 1, 
/* out0348_had-eta8-phi17*/	3, 22, 2, 7, 38, 0, 5, 39, 1, 8, 
/* out0349_had-eta9-phi17*/	3, 38, 0, 7, 38, 1, 8, 38, 2, 1, 
/* out0350_had-eta10-phi17*/	2, 37, 0, 8, 38, 1, 6, 
/* out0351_had-eta11-phi17*/	5, 37, 0, 3, 37, 1, 3, 37, 2, 5, 107, 0, 13, 107, 1, 1, 
/* out0352_had-eta12-phi17*/	6, 36, 0, 2, 37, 1, 4, 37, 2, 2, 105, 0, 10, 105, 2, 2, 107, 0, 1, 
/* out0353_had-eta13-phi17*/	4, 36, 0, 2, 36, 2, 7, 105, 1, 6, 105, 2, 5, 
/* out0354_had-eta14-phi17*/	4, 36, 2, 6, 103, 0, 4, 103, 2, 2, 105, 1, 2, 
/* out0355_had-eta15-phi17*/	6, 35, 2, 1, 36, 1, 1, 36, 2, 1, 43, 0, 2, 43, 1, 2, 103, 2, 7, 
/* out0356_had-eta16-phi17*/	5, 35, 2, 3, 43, 1, 2, 103, 1, 1, 103, 2, 4, 108, 0, 2, 
/* out0357_had-eta17-phi17*/	5, 35, 2, 2, 42, 0, 2, 102, 2, 2, 108, 0, 1, 108, 1, 3, 
/* out0358_had-eta18-phi17*/	3, 42, 0, 3, 102, 2, 4, 108, 1, 1, 
/* out0359_had-eta19-phi17*/	1, 42, 0, 1, 
/* out0360_had-eta0-phi18*/	0, 
/* out0361_had-eta1-phi18*/	1, 147, 0, 1, 
/* out0362_had-eta2-phi18*/	2, 146, 0, 1, 147, 0, 7, 
/* out0363_had-eta3-phi18*/	1, 146, 0, 4, 
/* out0364_had-eta4-phi18*/	1, 146, 0, 3, 
/* out0365_had-eta5-phi18*/	4, 24, 0, 3, 24, 1, 6, 28, 0, 7, 28, 2, 8, 
/* out0366_had-eta6-phi18*/	7, 23, 0, 10, 23, 1, 5, 24, 1, 1, 26, 0, 1, 26, 2, 2, 28, 1, 2, 28, 2, 8, 
/* out0367_had-eta7-phi18*/	3, 22, 0, 9, 23, 1, 9, 26, 2, 5, 
/* out0368_had-eta8-phi18*/	3, 22, 0, 4, 22, 1, 9, 22, 2, 7, 
/* out0369_had-eta9-phi18*/	6, 21, 0, 6, 21, 2, 6, 22, 1, 2, 22, 2, 1, 38, 0, 1, 38, 1, 1, 
/* out0370_had-eta10-phi18*/	4, 21, 1, 1, 21, 2, 10, 37, 0, 3, 106, 0, 1, 
/* out0371_had-eta11-phi18*/	6, 20, 2, 3, 37, 0, 2, 37, 1, 6, 106, 0, 6, 106, 2, 11, 107, 0, 1, 
/* out0372_had-eta12-phi18*/	7, 20, 2, 2, 36, 0, 4, 37, 1, 3, 105, 0, 5, 105, 1, 1, 106, 1, 1, 106, 2, 5, 
/* out0373_had-eta13-phi18*/	4, 36, 0, 6, 36, 1, 2, 104, 2, 4, 105, 1, 7, 
/* out0374_had-eta14-phi18*/	3, 36, 1, 6, 103, 0, 8, 104, 2, 1, 
/* out0375_had-eta15-phi18*/	5, 35, 0, 4, 36, 1, 1, 103, 0, 2, 103, 1, 4, 103, 2, 1, 
/* out0376_had-eta16-phi18*/	4, 35, 0, 1, 35, 2, 4, 102, 0, 1, 103, 1, 5, 
/* out0377_had-eta17-phi18*/	3, 35, 2, 4, 102, 0, 4, 102, 2, 2, 
/* out0378_had-eta18-phi18*/	3, 35, 2, 2, 42, 0, 1, 102, 2, 6, 
/* out0379_had-eta19-phi18*/	1, 102, 2, 1, 
/* out0380_had-eta0-phi19*/	0, 
/* out0381_had-eta1-phi19*/	1, 149, 0, 1, 
/* out0382_had-eta2-phi19*/	2, 148, 0, 1, 149, 0, 7, 
/* out0383_had-eta3-phi19*/	1, 148, 0, 4, 
/* out0384_had-eta4-phi19*/	1, 148, 0, 3, 
/* out0385_had-eta5-phi19*/	4, 27, 0, 2, 27, 2, 3, 28, 0, 9, 28, 1, 5, 
/* out0386_had-eta6-phi19*/	3, 26, 0, 13, 27, 2, 6, 28, 1, 9, 
/* out0387_had-eta7-phi19*/	5, 22, 0, 1, 25, 0, 2, 26, 0, 1, 26, 1, 11, 26, 2, 9, 
/* out0388_had-eta8-phi19*/	4, 22, 0, 1, 22, 1, 5, 25, 0, 4, 25, 2, 11, 
/* out0389_had-eta9-phi19*/	3, 21, 0, 10, 21, 1, 3, 25, 2, 4, 
/* out0390_had-eta10-phi19*/	2, 20, 0, 2, 21, 1, 12, 
/* out0391_had-eta11-phi19*/	4, 20, 0, 7, 20, 2, 4, 106, 0, 9, 106, 1, 9, 
/* out0392_had-eta12-phi19*/	4, 20, 1, 2, 20, 2, 7, 104, 0, 7, 106, 1, 6, 
/* out0393_had-eta13-phi19*/	7, 14, 2, 1, 20, 1, 1, 36, 0, 2, 36, 1, 3, 104, 0, 3, 104, 1, 1, 104, 2, 7, 
/* out0394_had-eta14-phi19*/	5, 14, 2, 3, 36, 1, 3, 103, 0, 2, 104, 1, 2, 104, 2, 4, 
/* out0395_had-eta15-phi19*/	3, 35, 0, 5, 98, 2, 3, 103, 1, 4, 
/* out0396_had-eta16-phi19*/	5, 35, 0, 3, 35, 1, 2, 98, 2, 2, 102, 0, 2, 103, 1, 2, 
/* out0397_had-eta17-phi19*/	2, 35, 1, 4, 102, 0, 5, 
/* out0398_had-eta18-phi19*/	4, 35, 1, 2, 102, 0, 1, 102, 1, 4, 102, 2, 1, 
/* out0399_had-eta19-phi19*/	1, 102, 1, 2, 
/* out0400_had-eta0-phi20*/	0, 
/* out0401_had-eta1-phi20*/	1, 149, 0, 1, 
/* out0402_had-eta2-phi20*/	2, 148, 0, 1, 149, 0, 7, 
/* out0403_had-eta3-phi20*/	1, 148, 0, 4, 
/* out0404_had-eta4-phi20*/	1, 148, 0, 3, 
/* out0405_had-eta5-phi20*/	3, 27, 0, 14, 27, 1, 3, 27, 2, 1, 
/* out0406_had-eta6-phi20*/	6, 26, 0, 1, 26, 1, 1, 27, 1, 13, 27, 2, 6, 33, 0, 6, 33, 2, 1, 
/* out0407_had-eta7-phi20*/	4, 25, 0, 3, 26, 1, 4, 33, 0, 1, 33, 2, 15, 
/* out0408_had-eta8-phi20*/	3, 25, 0, 7, 25, 1, 11, 25, 2, 1, 
/* out0409_had-eta9-phi20*/	3, 25, 1, 5, 29, 0, 7, 29, 2, 2, 
/* out0410_had-eta10-phi20*/	2, 20, 0, 1, 29, 2, 12, 
/* out0411_had-eta11-phi20*/	5, 20, 0, 6, 20, 1, 5, 29, 2, 1, 101, 0, 8, 101, 2, 8, 
/* out0412_had-eta12-phi20*/	4, 14, 0, 1, 20, 1, 8, 101, 2, 8, 104, 0, 4, 
/* out0413_had-eta13-phi20*/	4, 14, 0, 6, 14, 2, 2, 104, 0, 2, 104, 1, 8, 
/* out0414_had-eta14-phi20*/	3, 14, 2, 7, 98, 0, 4, 104, 1, 5, 
/* out0415_had-eta15-phi20*/	4, 14, 2, 3, 35, 0, 2, 98, 0, 3, 98, 2, 4, 
/* out0416_had-eta16-phi20*/	3, 35, 0, 1, 35, 1, 4, 98, 2, 6, 
/* out0417_had-eta17-phi20*/	4, 35, 1, 4, 98, 2, 1, 102, 0, 3, 102, 1, 2, 
/* out0418_had-eta18-phi20*/	1, 102, 1, 6, 
/* out0419_had-eta19-phi20*/	1, 102, 1, 2, 
/* out0420_had-eta0-phi21*/	0, 
/* out0421_had-eta1-phi21*/	1, 151, 0, 1, 
/* out0422_had-eta2-phi21*/	2, 150, 0, 1, 151, 0, 7, 
/* out0423_had-eta3-phi21*/	1, 150, 0, 4, 
/* out0424_had-eta4-phi21*/	1, 150, 0, 3, 
/* out0425_had-eta5-phi21*/	3, 34, 0, 14, 34, 1, 1, 34, 2, 3, 
/* out0426_had-eta6-phi21*/	6, 31, 0, 1, 31, 2, 1, 33, 0, 7, 33, 1, 1, 34, 1, 6, 34, 2, 13, 
/* out0427_had-eta7-phi21*/	4, 30, 0, 3, 31, 2, 4, 33, 0, 2, 33, 1, 15, 
/* out0428_had-eta8-phi21*/	3, 30, 0, 7, 30, 1, 1, 30, 2, 11, 
/* out0429_had-eta9-phi21*/	3, 29, 0, 8, 29, 1, 2, 30, 2, 5, 
/* out0430_had-eta10-phi21*/	4, 15, 0, 1, 29, 0, 1, 29, 1, 13, 29, 2, 1, 
/* out0431_had-eta11-phi21*/	5, 15, 0, 6, 15, 2, 5, 29, 1, 1, 101, 0, 8, 101, 1, 8, 
/* out0432_had-eta12-phi21*/	4, 14, 0, 1, 15, 2, 8, 99, 0, 4, 101, 1, 8, 
/* out0433_had-eta13-phi21*/	4, 14, 0, 7, 14, 1, 1, 99, 0, 2, 99, 2, 8, 
/* out0434_had-eta14-phi21*/	3, 14, 1, 7, 98, 0, 4, 99, 2, 5, 
/* out0435_had-eta15-phi21*/	4, 7, 0, 2, 14, 1, 3, 98, 0, 4, 98, 1, 4, 
/* out0436_had-eta16-phi21*/	3, 7, 0, 1, 7, 2, 4, 98, 1, 6, 
/* out0437_had-eta17-phi21*/	4, 7, 2, 4, 98, 1, 1, 128, 0, 3, 128, 2, 2, 
/* out0438_had-eta18-phi21*/	1, 128, 2, 6, 
/* out0439_had-eta19-phi21*/	1, 128, 2, 2, 
/* out0440_had-eta0-phi22*/	0, 
/* out0441_had-eta1-phi22*/	1, 151, 0, 1, 
/* out0442_had-eta2-phi22*/	2, 150, 0, 1, 151, 0, 7, 
/* out0443_had-eta3-phi22*/	1, 150, 0, 4, 
/* out0444_had-eta4-phi22*/	1, 150, 0, 3, 
/* out0445_had-eta5-phi22*/	4, 32, 0, 9, 32, 2, 5, 34, 0, 2, 34, 1, 3, 
/* out0446_had-eta6-phi22*/	3, 31, 0, 13, 32, 2, 9, 34, 1, 6, 
/* out0447_had-eta7-phi22*/	5, 17, 0, 1, 30, 0, 2, 31, 0, 1, 31, 1, 9, 31, 2, 11, 
/* out0448_had-eta8-phi22*/	4, 17, 0, 1, 17, 2, 5, 30, 0, 4, 30, 1, 11, 
/* out0449_had-eta9-phi22*/	3, 16, 0, 10, 16, 2, 3, 30, 1, 4, 
/* out0450_had-eta10-phi22*/	2, 15, 0, 2, 16, 2, 12, 
/* out0451_had-eta11-phi22*/	4, 15, 0, 7, 15, 1, 4, 100, 0, 9, 100, 2, 9, 
/* out0452_had-eta12-phi22*/	4, 15, 1, 7, 15, 2, 2, 99, 0, 7, 100, 2, 6, 
/* out0453_had-eta13-phi22*/	8, 8, 0, 2, 8, 2, 3, 14, 0, 1, 14, 1, 2, 15, 2, 1, 99, 0, 3, 99, 1, 7, 99, 2, 1, 
/* out0454_had-eta14-phi22*/	6, 8, 2, 3, 14, 1, 3, 98, 0, 1, 99, 1, 4, 99, 2, 2, 129, 0, 2, 
/* out0455_had-eta15-phi22*/	3, 7, 0, 5, 98, 1, 3, 129, 2, 4, 
/* out0456_had-eta16-phi22*/	5, 7, 0, 3, 7, 2, 2, 98, 1, 2, 128, 0, 2, 129, 2, 2, 
/* out0457_had-eta17-phi22*/	2, 7, 2, 4, 128, 0, 5, 
/* out0458_had-eta18-phi22*/	4, 7, 2, 2, 128, 0, 1, 128, 1, 1, 128, 2, 4, 
/* out0459_had-eta19-phi22*/	1, 128, 2, 2, 
/* out0460_had-eta0-phi23*/	0, 
/* out0461_had-eta1-phi23*/	1, 153, 0, 1, 
/* out0462_had-eta2-phi23*/	2, 152, 0, 1, 153, 0, 7, 
/* out0463_had-eta3-phi23*/	1, 152, 0, 4, 
/* out0464_had-eta4-phi23*/	1, 152, 0, 3, 
/* out0465_had-eta5-phi23*/	4, 19, 0, 3, 19, 2, 6, 32, 0, 7, 32, 1, 8, 
/* out0466_had-eta6-phi23*/	7, 18, 0, 10, 18, 2, 5, 19, 2, 1, 31, 0, 1, 31, 1, 2, 32, 1, 8, 32, 2, 2, 
/* out0467_had-eta7-phi23*/	3, 17, 0, 9, 18, 2, 9, 31, 1, 5, 
/* out0468_had-eta8-phi23*/	3, 17, 0, 4, 17, 1, 7, 17, 2, 9, 
/* out0469_had-eta9-phi23*/	6, 10, 0, 1, 10, 2, 1, 16, 0, 6, 16, 1, 6, 17, 1, 1, 17, 2, 2, 
/* out0470_had-eta10-phi23*/	4, 9, 0, 3, 16, 1, 10, 16, 2, 1, 100, 0, 1, 
/* out0471_had-eta11-phi23*/	6, 9, 0, 2, 9, 2, 6, 15, 1, 3, 100, 0, 6, 100, 1, 11, 131, 1, 1, 
/* out0472_had-eta12-phi23*/	7, 8, 0, 4, 9, 2, 3, 15, 1, 2, 100, 1, 5, 100, 2, 1, 130, 0, 5, 130, 2, 1, 
/* out0473_had-eta13-phi23*/	4, 8, 0, 6, 8, 2, 2, 99, 1, 4, 130, 2, 7, 
/* out0474_had-eta14-phi23*/	3, 8, 2, 6, 99, 1, 1, 129, 0, 8, 
/* out0475_had-eta15-phi23*/	5, 7, 0, 4, 8, 2, 1, 129, 0, 2, 129, 1, 1, 129, 2, 4, 
/* out0476_had-eta16-phi23*/	4, 7, 0, 1, 7, 1, 4, 128, 0, 1, 129, 2, 5, 
/* out0477_had-eta17-phi23*/	3, 7, 1, 4, 128, 0, 4, 128, 1, 2, 
/* out0478_had-eta18-phi23*/	3, 0, 0, 1, 7, 1, 2, 128, 1, 6, 
/* out0479_had-eta19-phi23*/	1, 128, 1, 1, 
};