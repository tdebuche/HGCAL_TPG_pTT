parameter integer matrixH [0:7586] = {
/* num inputs = 116(in0-in115) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 13 */
//* total number of input in adders 2368 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	0,
/* out0003_em-eta3-phi0*/	0,
/* out0004_em-eta4-phi0*/	0,
/* out0005_em-eta5-phi0*/	3,75,1,1,85,1,8,85,2,15,
/* out0006_em-eta6-phi0*/	3,75,0,14,75,1,7,75,2,3,
/* out0007_em-eta7-phi0*/	8,54,0,1,54,1,3,63,1,6,63,2,14,65,0,6,65,1,6,75,0,2,75,2,4,
/* out0008_em-eta8-phi0*/	6,54,0,14,54,1,3,54,2,2,54,1,1,65,0,10,65,2,4,
/* out0009_em-eta9-phi0*/	6,45,0,5,45,1,3,54,0,1,54,2,2,54,0,11,54,1,2,
/* out0010_em-eta10-phi0*/	6,45,0,11,45,2,1,43,0,1,43,1,1,54,0,5,54,2,2,
/* out0011_em-eta11-phi0*/	6,35,0,4,35,1,2,45,2,1,104,0,11,104,1,1,43,0,8,
/* out0012_em-eta12-phi0*/	6,35,0,9,104,0,2,104,1,2,104,2,9,43,0,5,43,2,1,
/* out0013_em-eta13-phi0*/	7,25,0,1,25,1,1,35,0,1,35,2,1,96,0,8,104,2,3,32,0,3,
/* out0014_em-eta14-phi0*/	5,25,0,6,96,0,4,96,1,1,96,2,5,32,0,6,
/* out0015_em-eta15-phi0*/	4,25,0,4,88,0,2,96,2,6,32,0,2,
/* out0016_em-eta16-phi0*/	3,17,2,1,88,0,7,22,0,2,
/* out0017_em-eta17-phi0*/	5,17,0,1,17,2,4,88,0,2,88,2,4,22,0,3,
/* out0018_em-eta18-phi0*/	2,88,2,5,22,0,1,
/* out0019_em-eta19-phi0*/	1,88,2,1,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	0,
/* out0023_em-eta3-phi1*/	0,
/* out0024_em-eta4-phi1*/	0,
/* out0025_em-eta5-phi1*/	5,85,1,8,85,2,1,86,0,11,86,1,7,86,2,1,
/* out0026_em-eta6-phi1*/	7,64,1,1,75,1,8,75,2,6,76,0,4,76,1,2,86,0,5,86,2,4,
/* out0027_em-eta7-phi1*/	8,54,1,3,63,1,10,63,2,2,64,0,12,64,1,1,65,1,10,75,2,3,76,0,11,
/* out0028_em-eta8-phi1*/	7,54,1,7,54,2,9,55,0,3,64,0,2,54,1,2,65,2,12,66,0,6,
/* out0029_em-eta9-phi1*/	6,45,1,11,54,2,3,55,0,5,54,1,11,54,2,4,66,0,1,
/* out0030_em-eta10-phi1*/	6,45,1,2,45,2,12,46,0,1,43,1,4,54,2,9,55,0,1,
/* out0031_em-eta11-phi1*/	8,35,1,10,45,2,1,104,0,3,104,1,5,111,2,10,43,0,1,43,1,8,43,2,2,
/* out0032_em-eta12-phi1*/	9,35,0,2,35,1,1,35,2,7,104,1,8,104,2,3,105,0,5,32,1,1,43,0,1,43,2,8,
/* out0033_em-eta13-phi1*/	9,25,1,5,35,2,3,96,0,4,96,1,4,104,2,1,105,0,1,105,2,3,32,0,1,32,1,7,
/* out0034_em-eta14-phi1*/	8,25,0,3,25,1,3,25,2,1,96,1,8,96,2,1,32,0,3,32,1,1,32,2,2,
/* out0035_em-eta15-phi1*/	10,25,0,2,25,2,4,88,0,2,88,1,1,96,1,2,96,2,4,97,0,1,22,1,1,32,0,1,32,2,4,
/* out0036_em-eta16-phi1*/	6,17,2,5,25,2,1,88,0,2,88,1,4,22,0,2,22,1,3,
/* out0037_em-eta17-phi1*/	6,17,0,3,17,2,3,88,0,1,88,1,4,88,2,1,22,0,4,
/* out0038_em-eta18-phi1*/	4,88,1,1,88,2,4,22,0,3,22,2,1,
/* out0039_em-eta19-phi1*/	2,22,0,1,22,2,1,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	0,
/* out0043_em-eta3-phi2*/	0,
/* out0044_em-eta4-phi2*/	0,
/* out0045_em-eta5-phi2*/	7,86,1,9,86,2,5,87,0,2,87,1,2,94,0,14,94,1,13,94,2,12,
/* out0046_em-eta6-phi2*/	7,64,1,3,71,0,4,71,1,2,71,2,2,76,1,12,86,2,6,87,0,10,
/* out0047_em-eta7-phi2*/	12,64,0,2,64,1,11,64,2,11,65,0,1,71,0,5,71,1,5,71,2,1,66,1,3,76,0,1,76,1,2,76,2,16,77,0,3,
/* out0048_em-eta8-phi2*/	7,55,0,2,55,1,13,64,2,5,65,0,1,66,0,6,66,1,10,66,2,4,
/* out0049_em-eta9-phi2*/	8,46,1,1,55,0,6,55,2,10,54,2,1,55,0,2,55,1,5,66,0,3,66,2,6,
/* out0050_em-eta10-phi2*/	7,45,2,1,46,0,8,46,1,6,111,2,1,55,0,11,55,1,2,55,2,1,
/* out0051_em-eta11-phi2*/	12,35,1,3,46,0,7,46,2,3,105,0,1,111,1,14,111,2,5,43,1,3,43,2,2,44,0,1,44,1,1,55,0,2,55,2,2,
/* out0052_em-eta12-phi2*/	7,35,2,4,36,0,5,36,1,1,105,0,9,105,1,3,43,2,3,44,0,7,
/* out0053_em-eta13-phi2*/	7,25,1,3,35,2,1,36,0,5,105,1,1,105,2,9,32,1,6,44,0,2,
/* out0054_em-eta14-phi2*/	7,25,1,4,25,2,3,96,1,1,97,0,6,105,2,2,32,1,1,32,2,6,
/* out0055_em-eta15-phi2*/	7,25,2,6,26,0,1,97,0,4,97,2,3,22,1,2,32,2,3,33,0,1,
/* out0056_em-eta16-phi2*/	5,17,0,3,17,2,3,88,1,2,97,2,4,22,1,5,
/* out0057_em-eta17-phi2*/	5,17,0,4,88,1,3,89,1,2,22,1,1,22,2,2,
/* out0058_em-eta18-phi2*/	4,88,1,1,88,2,1,89,1,2,22,2,3,
/* out0059_em-eta19-phi2*/	1,22,2,1,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	0,
/* out0063_em-eta3-phi3*/	0,
/* out0064_em-eta4-phi3*/	0,
/* out0065_em-eta5-phi3*/	7,87,1,11,94,0,2,94,1,3,94,2,4,95,0,16,95,1,4,95,2,8,
/* out0066_em-eta6-phi3*/	7,71,0,1,72,0,4,77,1,5,87,0,4,87,1,3,87,2,16,88,0,3,
/* out0067_em-eta7-phi3*/	11,65,0,6,65,1,13,65,2,1,71,0,6,71,1,9,71,2,13,72,0,3,72,2,1,77,0,11,77,1,8,77,2,5,
/* out0068_em-eta8-phi3*/	11,55,1,3,55,2,1,56,1,3,65,0,8,65,2,7,66,1,3,66,2,4,67,0,5,67,1,4,77,0,2,77,2,3,
/* out0069_em-eta9-phi3*/	7,46,1,1,55,2,5,56,0,11,56,1,1,55,1,5,66,2,2,67,0,9,
/* out0070_em-eta10-phi3*/	9,46,1,8,46,2,4,56,0,2,111,1,1,112,0,1,112,1,1,55,1,4,55,2,9,56,0,1,
/* out0071_em-eta11-phi3*/	10,36,1,3,46,2,9,47,0,1,111,1,1,112,0,15,112,1,3,112,2,5,44,1,7,55,2,4,56,0,1,
/* out0072_em-eta12-phi3*/	9,36,0,2,36,1,8,36,2,1,105,1,7,106,0,1,112,2,5,44,0,4,44,1,3,44,2,3,
/* out0073_em-eta13-phi3*/	9,36,0,4,36,2,5,105,1,5,105,2,2,106,0,3,106,2,1,33,1,1,44,0,2,44,2,4,
/* out0074_em-eta14-phi3*/	9,25,2,1,26,0,2,26,1,3,36,2,1,97,0,4,97,1,5,32,2,1,33,0,5,33,1,2,
/* out0075_em-eta15-phi3*/	5,26,0,6,97,0,1,97,1,4,97,2,3,33,0,5,
/* out0076_em-eta16-phi3*/	6,17,0,2,26,0,3,89,2,1,97,2,5,22,1,3,33,0,1,
/* out0077_em-eta17-phi3*/	5,17,0,3,89,1,2,89,2,3,22,1,1,22,2,4,
/* out0078_em-eta18-phi3*/	2,89,1,4,22,2,3,
/* out0079_em-eta19-phi3*/	2,89,1,1,22,2,1,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	0,
/* out0083_em-eta3-phi4*/	0,
/* out0084_em-eta4-phi4*/	0,
/* out0085_em-eta5-phi4*/	6,88,1,6,95,1,12,95,2,8,96,0,13,96,1,1,96,2,2,
/* out0086_em-eta6-phi4*/	5,72,0,2,72,1,6,88,0,12,88,1,8,88,2,8,
/* out0087_em-eta7-phi4*/	13,65,1,3,65,2,3,66,0,2,66,1,4,72,0,7,72,1,6,72,2,14,77,1,3,77,2,7,78,0,8,78,1,4,88,0,1,88,2,2,
/* out0088_em-eta8-phi4*/	7,56,1,6,65,2,5,66,0,10,67,1,12,67,2,2,77,2,1,78,0,5,
/* out0089_em-eta9-phi4*/	6,56,0,2,56,1,6,56,2,10,56,1,2,67,0,2,67,2,12,
/* out0090_em-eta10-phi4*/	6,47,0,2,47,1,7,56,0,1,56,2,4,56,0,7,56,1,6,
/* out0091_em-eta11-phi4*/	8,47,0,11,47,1,1,47,2,1,112,1,11,112,2,1,44,1,3,56,0,7,56,2,1,
/* out0092_em-eta12-phi4*/	12,36,1,4,36,2,3,37,0,1,47,0,2,47,2,1,106,0,7,106,1,1,112,1,1,112,2,5,44,1,2,44,2,6,45,0,2,
/* out0093_em-eta13-phi4*/	8,36,2,6,37,0,2,106,0,5,106,1,1,106,2,4,33,1,3,44,2,3,45,0,1,
/* out0094_em-eta14-phi4*/	6,26,1,7,97,1,2,98,0,1,106,2,5,33,0,1,33,1,6,
/* out0095_em-eta15-phi4*/	7,26,0,2,26,1,2,26,2,2,97,1,4,98,0,3,33,0,2,33,2,3,
/* out0096_em-eta16-phi4*/	10,26,0,2,26,2,3,89,2,3,97,1,1,97,2,1,98,0,1,98,2,1,23,2,1,33,0,1,33,2,2,
/* out0097_em-eta17-phi4*/	2,89,2,6,23,1,3,
/* out0098_em-eta18-phi4*/	3,89,0,2,89,1,3,23,1,3,
/* out0099_em-eta19-phi4*/	1,89,1,1,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	0,
/* out0103_em-eta3-phi5*/	0,
/* out0104_em-eta4-phi5*/	0,
/* out0105_em-eta5-phi5*/	4,89,1,2,96,0,3,96,1,15,96,2,13,
/* out0106_em-eta6-phi5*/	8,72,1,1,73,0,1,73,1,2,88,1,2,88,2,6,89,0,14,89,1,6,96,2,1,
/* out0107_em-eta7-phi5*/	11,66,1,11,66,2,1,72,1,3,72,2,1,73,0,15,73,1,4,73,2,8,78,0,1,78,1,12,78,2,8,89,0,2,
/* out0108_em-eta8-phi5*/	9,57,1,3,66,0,4,66,1,1,66,2,15,67,2,1,68,0,2,68,1,7,78,0,2,78,2,8,
/* out0109_em-eta9-phi5*/	7,56,2,2,57,0,10,57,1,5,56,1,2,67,2,1,68,0,13,68,1,1,
/* out0110_em-eta10-phi5*/	6,47,1,8,47,2,1,57,0,6,56,1,6,56,2,7,68,0,1,
/* out0111_em-eta11-phi5*/	6,47,2,12,113,0,15,113,1,5,113,2,1,45,1,3,56,2,8,
/* out0112_em-eta12-phi5*/	8,37,0,2,37,1,8,47,2,1,106,1,5,113,0,1,113,2,7,45,0,5,45,1,5,
/* out0113_em-eta13-phi5*/	5,37,0,8,106,1,9,106,2,2,33,1,1,45,0,7,
/* out0114_em-eta14-phi5*/	8,26,1,4,26,2,1,37,0,3,98,0,5,106,2,4,33,1,3,33,2,3,45,0,1,
/* out0115_em-eta15-phi5*/	4,26,2,6,98,0,6,98,2,1,33,2,6,
/* out0116_em-eta16-phi5*/	4,26,2,4,98,2,5,23,2,4,33,2,2,
/* out0117_em-eta17-phi5*/	5,89,0,3,89,2,3,98,2,1,23,1,1,23,2,2,
/* out0118_em-eta18-phi5*/	2,89,0,10,23,1,3,
/* out0119_em-eta19-phi5*/	3,89,0,1,89,1,1,23,1,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	0,
/* out0123_em-eta3-phi6*/	0,
/* out0124_em-eta4-phi6*/	0,
/* out0125_em-eta5-phi6*/	4,89,1,2,97,0,16,97,1,11,97,2,13,
/* out0126_em-eta6-phi6*/	8,73,1,2,74,0,1,74,1,1,89,1,6,89,2,14,90,0,6,90,1,2,97,2,1,
/* out0127_em-eta7-phi6*/	10,67,0,1,67,1,11,73,1,8,73,2,8,74,0,10,74,2,1,79,0,8,79,1,12,79,2,1,89,2,2,
/* out0128_em-eta8-phi6*/	9,57,1,3,67,0,15,67,1,1,67,2,4,68,1,7,68,2,2,69,0,1,79,0,8,79,2,2,
/* out0129_em-eta9-phi6*/	7,57,1,5,57,2,10,58,0,2,57,1,2,68,1,1,68,2,13,69,0,1,
/* out0130_em-eta10-phi6*/	6,48,0,1,48,1,8,57,2,6,57,0,7,57,1,6,68,2,1,
/* out0131_em-eta11-phi6*/	6,48,0,12,113,1,11,113,2,1,114,0,1,45,1,3,57,0,8,
/* out0132_em-eta12-phi6*/	7,37,1,8,37,2,2,48,0,1,107,0,5,113,2,7,45,1,5,45,2,5,
/* out0133_em-eta13-phi6*/	5,37,2,8,107,0,9,107,2,2,34,1,1,45,2,7,
/* out0134_em-eta14-phi6*/	8,27,0,1,27,1,4,37,2,3,98,1,5,107,2,4,34,0,3,34,1,3,45,2,1,
/* out0135_em-eta15-phi6*/	4,27,0,6,98,1,6,98,2,1,34,0,6,
/* out0136_em-eta16-phi6*/	4,27,0,4,98,2,5,23,2,4,34,0,2,
/* out0137_em-eta17-phi6*/	5,90,1,1,90,2,3,98,2,1,23,0,2,23,2,3,
/* out0138_em-eta18-phi6*/	3,90,1,4,23,0,1,23,1,3,
/* out0139_em-eta19-phi6*/	2,90,1,2,23,1,1,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	0,
/* out0143_em-eta3-phi7*/	0,
/* out0144_em-eta4-phi7*/	0,
/* out0145_em-eta5-phi7*/	6,90,1,6,97,1,5,97,2,2,98,0,16,98,1,7,98,2,8,
/* out0146_em-eta6-phi7*/	4,74,1,7,90,0,8,90,1,8,90,2,12,
/* out0147_em-eta7-phi7*/	13,67,1,4,67,2,2,68,0,3,68,1,3,74,0,5,74,1,6,74,2,14,79,1,4,79,2,8,80,0,7,80,1,3,90,0,2,90,2,1,
/* out0148_em-eta8-phi7*/	7,58,1,6,67,2,10,68,0,5,69,0,2,69,1,12,79,2,5,80,0,1,
/* out0149_em-eta9-phi7*/	6,58,0,10,58,1,6,58,2,2,57,1,2,69,0,12,69,2,2,
/* out0150_em-eta10-phi7*/	6,48,1,7,48,2,2,58,0,4,58,2,1,57,1,6,57,2,7,
/* out0151_em-eta11-phi7*/	9,48,0,1,48,1,1,48,2,11,114,0,14,114,1,5,114,2,2,46,1,3,57,0,1,57,2,7,
/* out0152_em-eta12-phi7*/	12,37,2,1,38,0,3,38,1,4,48,0,1,48,2,2,107,0,1,107,1,7,114,0,1,114,2,5,45,2,2,46,0,6,46,1,2,
/* out0153_em-eta13-phi7*/	8,37,2,2,38,0,6,107,0,1,107,1,5,107,2,4,34,1,3,45,2,1,46,0,3,
/* out0154_em-eta14-phi7*/	6,27,1,7,98,1,1,99,0,2,107,2,5,34,1,6,34,2,1,
/* out0155_em-eta15-phi7*/	7,27,0,2,27,1,2,27,2,2,98,1,3,99,0,4,34,0,3,34,2,2,
/* out0156_em-eta16-phi7*/	10,27,0,3,27,2,2,90,2,3,98,1,1,98,2,1,99,0,1,99,2,1,23,2,1,34,0,2,34,2,1,
/* out0157_em-eta17-phi7*/	3,90,2,5,23,0,7,23,2,1,
/* out0158_em-eta18-phi7*/	3,90,1,4,23,0,5,23,1,1,
/* out0159_em-eta19-phi7*/	1,90,1,1,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	0,
/* out0163_em-eta3-phi8*/	0,
/* out0164_em-eta4-phi8*/	0,
/* out0165_em-eta5-phi8*/	6,91,1,11,98,1,9,98,2,8,99,0,4,99,1,3,99,2,2,
/* out0166_em-eta6-phi8*/	7,74,1,1,75,2,1,80,1,5,90,2,3,91,0,16,91,1,3,91,2,4,
/* out0167_em-eta7-phi8*/	11,68,0,1,68,1,13,68,2,6,74,1,1,74,2,1,75,0,13,75,1,9,75,2,6,80,0,5,80,1,8,80,2,11,
/* out0168_em-eta8-phi8*/	11,58,1,3,59,0,1,59,1,3,68,0,7,68,2,8,69,1,4,69,2,5,70,0,4,70,1,3,80,0,3,80,2,2,
/* out0169_em-eta9-phi8*/	7,49,1,1,58,1,1,58,2,11,59,0,5,58,1,5,69,2,9,70,0,2,
/* out0170_em-eta10-phi8*/	8,49,0,4,49,1,8,58,2,2,114,1,2,115,0,1,57,2,1,58,0,9,58,1,4,
/* out0171_em-eta11-phi8*/	9,38,1,3,48,2,1,49,0,9,114,1,9,114,2,4,115,0,1,46,1,7,57,2,1,58,0,4,
/* out0172_em-eta12-phi8*/	9,38,0,1,38,1,8,38,2,2,107,1,1,108,0,7,114,2,5,46,0,3,46,1,3,46,2,4,
/* out0173_em-eta13-phi8*/	9,38,0,5,38,2,4,107,1,3,107,2,1,108,0,5,108,2,2,34,1,1,46,0,4,46,2,2,
/* out0174_em-eta14-phi8*/	9,27,1,3,27,2,2,28,0,1,38,0,1,99,0,5,99,1,4,34,1,2,34,2,5,35,0,1,
/* out0175_em-eta15-phi8*/	5,27,2,6,99,0,4,99,1,1,99,2,2,34,2,5,
/* out0176_em-eta16-phi8*/	6,18,1,2,27,2,3,90,2,1,99,2,5,24,1,3,34,2,1,
/* out0177_em-eta17-phi8*/	5,18,1,3,90,0,4,90,2,4,24,0,4,24,1,1,
/* out0178_em-eta18-phi8*/	4,90,0,3,90,1,2,23,0,1,24,0,3,
/* out0179_em-eta19-phi8*/	2,90,1,1,24,0,1,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	0,
/* out0183_em-eta3-phi9*/	0,
/* out0184_em-eta4-phi9*/	0,
/* out0185_em-eta5-phi9*/	7,91,1,2,91,2,2,92,0,5,92,1,9,99,0,12,99,1,13,99,2,14,
/* out0186_em-eta6-phi9*/	7,69,1,3,75,0,2,75,1,2,75,2,4,81,1,12,91,2,10,92,0,6,
/* out0187_em-eta7-phi9*/	12,68,2,1,69,0,11,69,1,11,69,2,2,75,0,1,75,1,5,75,2,5,70,1,3,80,2,3,81,0,16,81,1,2,81,2,1,
/* out0188_em-eta8-phi9*/	7,59,1,13,59,2,2,68,2,1,69,0,5,70,0,4,70,1,10,70,2,6,
/* out0189_em-eta9-phi9*/	8,49,1,1,59,0,10,59,2,6,58,1,5,58,2,2,59,0,1,70,0,6,70,2,3,
/* out0190_em-eta10-phi9*/	7,49,1,6,49,2,8,50,0,1,115,0,1,58,0,1,58,1,2,58,2,11,
/* out0191_em-eta11-phi9*/	12,39,1,3,49,0,3,49,2,7,108,1,1,115,0,11,115,2,8,46,1,1,46,2,1,47,0,2,47,1,3,58,0,2,58,2,2,
/* out0192_em-eta12-phi9*/	7,38,1,1,38,2,5,39,0,4,108,0,3,108,1,9,46,2,7,47,0,3,
/* out0193_em-eta13-phi9*/	7,28,1,3,38,2,5,39,0,1,108,0,1,108,2,9,35,1,6,46,2,2,
/* out0194_em-eta14-phi9*/	7,28,0,3,28,1,4,99,1,6,100,0,1,108,2,2,35,0,6,35,1,1,
/* out0195_em-eta15-phi9*/	7,27,2,1,28,0,6,99,1,4,99,2,3,24,1,2,34,2,1,35,0,3,
/* out0196_em-eta16-phi9*/	5,18,1,3,18,2,3,91,0,2,99,2,4,24,1,5,
/* out0197_em-eta17-phi9*/	5,18,1,4,90,0,4,91,0,3,24,0,2,24,1,1,
/* out0198_em-eta18-phi9*/	4,90,0,5,90,1,1,91,0,1,24,0,3,
/* out0199_em-eta19-phi9*/	1,24,0,1,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	0,
/* out0203_em-eta3-phi10*/	0,
/* out0204_em-eta4-phi10*/	0,
/* out0205_em-eta5-phi10*/	5,92,0,1,92,1,7,92,2,11,93,0,8,93,2,1,
/* out0206_em-eta6-phi10*/	8,69,1,1,70,0,1,81,1,2,81,2,4,82,0,6,82,1,8,92,0,4,92,2,5,
/* out0207_em-eta7-phi10*/	8,60,1,3,69,1,1,69,2,12,70,0,10,70,2,2,71,1,10,81,2,11,82,0,3,
/* out0208_em-eta8-phi10*/	7,59,2,3,60,0,9,60,1,7,69,2,2,59,1,2,70,2,6,71,0,12,
/* out0209_em-eta9-phi10*/	6,50,1,11,59,2,5,60,0,3,59,0,4,59,1,11,70,2,1,
/* out0210_em-eta10-phi10*/	6,49,2,1,50,0,12,50,1,2,47,1,4,58,2,1,59,0,9,
/* out0211_em-eta11-phi10*/	8,39,1,10,50,0,1,109,0,5,115,0,2,115,2,8,47,0,2,47,1,8,47,2,1,
/* out0212_em-eta12-phi10*/	8,39,0,7,39,1,1,39,2,2,108,1,5,109,0,8,35,1,1,47,0,8,47,2,1,
/* out0213_em-eta13-phi10*/	9,28,1,5,39,0,3,100,0,4,100,1,1,108,1,1,108,2,3,109,2,1,35,1,7,35,2,1,
/* out0214_em-eta14-phi10*/	7,28,0,1,28,1,3,28,2,3,100,0,8,35,0,2,35,1,1,35,2,3,
/* out0215_em-eta15-phi10*/	11,28,0,4,28,2,2,91,0,1,91,1,1,99,1,1,99,2,1,100,0,2,100,2,2,24,1,1,35,0,4,35,2,1,
/* out0216_em-eta16-phi10*/	6,18,2,5,28,0,1,91,0,4,91,1,2,24,1,3,24,2,2,
/* out0217_em-eta17-phi10*/	5,18,1,3,18,2,3,91,0,4,91,2,1,24,2,4,
/* out0218_em-eta18-phi10*/	4,91,0,1,91,2,3,24,0,1,24,2,3,
/* out0219_em-eta19-phi10*/	2,24,0,1,24,2,1,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	0,
/* out0223_em-eta3-phi11*/	0,
/* out0224_em-eta4-phi11*/	0,
/* out0225_em-eta5-phi11*/	4,82,1,1,83,1,4,93,0,8,93,2,15,
/* out0226_em-eta6-phi11*/	5,72,1,1,82,0,3,82,1,7,82,2,14,83,0,4,
/* out0227_em-eta7-phi11*/	12,60,1,3,60,2,1,61,0,2,61,1,4,70,0,5,70,2,14,71,1,6,71,2,6,72,0,4,72,1,3,82,0,4,82,2,2,
/* out0228_em-eta8-phi11*/	10,51,1,1,60,0,2,60,1,3,60,2,14,61,0,2,59,1,1,60,0,1,60,1,4,71,0,4,71,2,10,
/* out0229_em-eta9-phi11*/	9,50,1,3,50,2,5,51,0,4,51,1,3,60,0,2,60,2,1,59,1,2,59,2,11,60,0,3,
/* out0230_em-eta10-phi11*/	9,40,1,3,50,0,1,50,2,11,47,1,1,47,2,1,48,0,1,48,1,4,59,0,2,59,2,5,
/* out0231_em-eta11-phi11*/	9,39,1,2,39,2,5,40,0,4,40,1,1,50,0,1,109,0,1,109,1,10,47,2,8,48,0,3,
/* out0232_em-eta12-phi11*/	8,29,1,2,39,2,8,109,0,2,109,1,2,109,2,8,36,1,4,47,0,1,47,2,5,
/* out0233_em-eta13-phi11*/	10,28,1,1,28,2,1,29,0,3,29,1,2,39,0,1,39,2,1,100,1,7,109,2,3,35,2,3,36,0,4,
/* out0234_em-eta14-phi11*/	7,28,2,6,29,0,1,100,0,1,100,1,4,100,2,4,25,1,1,35,2,6,
/* out0235_em-eta15-phi11*/	7,19,1,3,28,2,4,91,1,1,100,2,6,25,0,1,25,1,3,35,2,2,
/* out0236_em-eta16-phi11*/	6,18,2,1,19,0,3,19,1,1,91,1,6,24,2,2,25,0,3,
/* out0237_em-eta17-phi11*/	6,18,1,1,18,2,4,19,0,1,91,1,2,91,2,4,24,2,3,
/* out0238_em-eta18-phi11*/	3,91,2,4,14,1,2,24,2,1,
/* out0239_em-eta19-phi11*/	1,14,1,3,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	0,
/* out0243_em-eta3-phi12*/	0,
/* out0244_em-eta4-phi12*/	0,
/* out0245_em-eta5-phi12*/	3,83,1,12,83,2,8,84,0,3,
/* out0246_em-eta6-phi12*/	6,72,1,7,72,2,3,73,0,1,73,1,1,83,0,12,83,2,6,
/* out0247_em-eta7-phi12*/	7,61,0,3,61,1,12,61,2,9,62,0,1,72,0,10,72,1,5,72,2,9,
/* out0248_em-eta8-phi12*/	8,51,1,8,51,2,2,61,0,9,61,2,2,60,0,1,60,1,12,60,2,5,72,0,2,
/* out0249_em-eta9-phi12*/	6,51,0,8,51,1,4,51,2,6,48,1,3,60,0,11,60,2,2,
/* out0250_em-eta10-phi12*/	6,40,1,10,40,2,1,51,0,4,48,0,2,48,1,9,48,2,3,
/* out0251_em-eta11-phi12*/	9,40,0,8,40,1,2,40,2,2,109,1,3,110,0,11,110,2,1,36,1,2,48,0,9,48,2,1,
/* out0252_em-eta12-phi12*/	10,29,1,7,40,0,3,101,0,5,101,1,2,109,1,1,109,2,4,110,0,1,110,2,1,36,1,9,36,2,1,
/* out0253_em-eta13-phi12*/	7,29,0,4,29,1,4,29,2,1,100,1,2,101,0,8,36,0,7,36,2,1,
/* out0254_em-eta14-phi12*/	10,19,1,1,29,0,6,92,0,1,92,1,1,100,1,2,100,2,3,101,0,1,101,2,1,25,1,4,36,0,3,
/* out0255_em-eta15-phi12*/	5,19,1,6,92,0,6,100,2,1,25,0,1,25,1,5,
/* out0256_em-eta16-phi12*/	5,19,0,4,19,1,2,91,1,3,92,0,4,25,0,5,
/* out0257_em-eta17-phi12*/	6,19,0,4,83,1,1,91,1,1,91,2,3,14,2,2,25,0,2,
/* out0258_em-eta18-phi12*/	4,83,1,4,91,2,1,14,1,3,14,2,1,
/* out0259_em-eta19-phi12*/	1,14,1,3,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	0,
/* out0263_em-eta3-phi13*/	0,
/* out0264_em-eta4-phi13*/	0,
/* out0265_em-eta5-phi13*/	6,73,1,3,73,2,1,74,0,1,83,2,1,84,0,13,84,2,14,
/* out0266_em-eta6-phi13*/	5,62,0,2,73,0,10,73,1,12,73,2,6,83,2,1,
/* out0267_em-eta7-phi13*/	8,52,1,7,61,2,4,62,0,12,62,2,9,61,1,15,61,2,1,72,2,4,73,0,5,
/* out0268_em-eta8-phi13*/	8,51,2,1,52,0,10,52,1,8,52,2,1,61,2,1,49,1,2,60,2,5,61,0,13,
/* out0269_em-eta9-phi13*/	6,41,1,9,51,2,7,52,0,3,49,0,4,49,1,9,60,2,4,
/* out0270_em-eta10-phi13*/	6,40,2,5,41,0,8,41,1,2,37,1,1,48,2,8,49,0,4,
/* out0271_em-eta11-phi13*/	10,30,1,5,40,2,8,102,0,1,110,0,4,110,2,12,36,1,1,37,0,2,37,1,5,48,0,1,48,2,4,
/* out0272_em-eta12-phi13*/	9,29,1,1,29,2,4,30,0,3,30,1,1,40,0,1,101,1,10,110,2,1,36,2,7,37,0,2,
/* out0273_em-eta13-phi13*/	7,29,2,8,101,0,2,101,1,1,101,2,7,26,1,1,36,0,1,36,2,7,
/* out0274_em-eta14-phi13*/	12,19,1,1,19,2,1,20,0,1,20,1,1,29,0,2,29,2,2,92,1,5,101,2,3,25,1,2,25,2,2,26,0,1,36,0,1,
/* out0275_em-eta15-phi13*/	7,19,1,2,19,2,4,92,0,3,92,1,3,92,2,1,25,1,1,25,2,5,
/* out0276_em-eta16-phi13*/	6,19,0,1,19,2,4,92,0,2,92,2,4,25,0,2,25,2,3,
/* out0277_em-eta17-phi13*/	7,19,0,3,19,2,1,83,1,2,83,2,4,92,2,1,14,2,3,25,0,2,
/* out0278_em-eta18-phi13*/	2,83,1,5,14,2,4,
/* out0279_em-eta19-phi13*/	1,14,1,2,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	0,
/* out0283_em-eta3-phi14*/	0,
/* out0284_em-eta4-phi14*/	0,
/* out0285_em-eta5-phi14*/	4,74,0,15,74,1,10,74,2,7,84,2,2,
/* out0286_em-eta6-phi14*/	7,53,0,2,53,1,1,62,0,1,62,2,1,62,1,12,73,2,9,74,2,8,
/* out0287_em-eta7-phi14*/	11,52,1,1,52,2,3,53,0,14,53,1,3,53,2,9,62,2,6,50,1,1,61,1,1,61,2,10,62,0,10,62,1,1,
/* out0288_em-eta8-phi14*/	10,42,1,6,52,0,2,52,2,12,53,2,1,49,1,2,49,2,1,50,0,3,50,1,5,61,0,3,61,2,5,
/* out0289_em-eta9-phi14*/	7,41,1,5,41,2,8,42,0,3,52,0,1,49,0,2,49,1,3,49,2,11,
/* out0290_em-eta10-phi14*/	8,30,1,1,41,0,8,41,2,6,102,1,1,37,1,5,37,2,1,49,0,6,49,2,2,
/* out0291_em-eta11-phi14*/	8,30,1,9,30,2,3,102,0,8,102,1,6,110,2,1,37,0,3,37,1,5,37,2,3,
/* out0292_em-eta12-phi14*/	7,30,0,9,30,2,1,101,1,3,102,0,7,102,2,3,26,1,2,37,0,7,
/* out0293_em-eta13-phi14*/	7,20,1,6,29,2,1,30,0,2,93,0,5,93,1,1,101,2,4,26,1,8,
/* out0294_em-eta14-phi14*/	7,20,0,3,20,1,4,92,1,3,93,0,5,101,2,1,26,0,6,26,1,1,
/* out0295_em-eta15-phi14*/	7,19,2,2,20,0,4,92,1,4,92,2,3,15,1,1,25,2,3,26,0,1,
/* out0296_em-eta16-phi14*/	6,11,1,2,19,2,3,84,0,1,92,2,6,15,1,2,25,2,2,
/* out0297_em-eta17-phi14*/	7,11,1,2,19,2,1,83,2,6,14,2,1,15,0,2,15,1,1,25,2,1,
/* out0298_em-eta18-phi14*/	3,83,1,3,83,2,2,14,2,4,
/* out0299_em-eta19-phi14*/	1,14,1,2,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	0,
/* out0303_em-eta3-phi15*/	0,
/* out0304_em-eta4-phi15*/	0,
/* out0305_em-eta5-phi15*/	2,63,1,13,74,1,5,
/* out0306_em-eta6-phi15*/	7,51,1,2,62,1,3,62,2,11,63,0,10,63,1,2,74,1,1,74,2,1,
/* out0307_em-eta7-phi15*/	10,43,0,1,43,1,5,53,1,12,53,2,5,50,1,5,50,2,3,51,0,2,51,1,3,62,0,6,62,2,5,
/* out0308_em-eta8-phi15*/	8,42,0,1,42,1,10,42,2,9,43,0,1,53,2,1,50,0,8,50,1,5,50,2,7,
/* out0309_em-eta9-phi15*/	7,31,1,5,41,2,1,42,0,11,42,2,1,38,1,10,49,2,2,50,0,5,
/* out0310_em-eta10-phi15*/	10,31,0,5,31,1,9,41,2,1,102,1,1,103,0,4,103,1,2,103,2,2,37,2,2,38,0,8,38,1,4,
/* out0311_em-eta11-phi15*/	11,21,1,1,30,2,7,31,0,4,102,1,8,102,2,5,103,0,6,103,1,5,103,2,1,27,1,2,37,2,8,38,0,1,
/* out0312_em-eta12-phi15*/	13,21,0,1,21,1,3,30,0,2,30,2,5,93,1,3,94,0,1,102,2,8,26,1,2,26,2,2,27,0,1,27,1,2,37,0,2,37,2,2,
/* out0313_em-eta13-phi15*/	7,20,1,4,20,2,5,93,0,2,93,1,8,93,2,1,26,1,2,26,2,5,
/* out0314_em-eta14-phi15*/	7,20,0,2,20,1,1,20,2,4,93,0,4,93,2,5,26,0,5,26,2,2,
/* out0315_em-eta15-phi15*/	8,11,2,1,20,0,5,84,0,2,84,1,3,92,2,1,93,2,1,15,1,4,26,0,2,
/* out0316_em-eta16-phi15*/	4,11,1,2,11,2,3,84,0,6,15,1,5,
/* out0317_em-eta17-phi15*/	4,11,1,4,83,2,2,84,0,3,15,0,3,
/* out0318_em-eta18-phi15*/	5,11,1,1,83,1,1,83,2,2,14,2,1,15,0,3,
/* out0319_em-eta19-phi15*/	1,14,1,1,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	0,
/* out0323_em-eta3-phi16*/	0,
/* out0324_em-eta4-phi16*/	0,
/* out0325_em-eta5-phi16*/	6,52,1,4,63,1,1,63,2,12,64,0,15,64,1,14,64,2,12,
/* out0326_em-eta6-phi16*/	11,43,1,1,43,2,1,44,0,3,44,1,2,44,2,1,51,1,7,51,2,5,52,0,3,52,1,4,63,0,6,63,2,4,
/* out0327_em-eta7-phi16*/	9,43,0,5,43,1,10,43,2,10,44,0,1,44,1,1,39,1,1,51,0,13,51,1,4,51,2,6,
/* out0328_em-eta8-phi16*/	6,32,1,9,42,2,4,43,0,9,39,0,2,39,1,12,50,2,6,
/* out0329_em-eta9-phi16*/	9,31,1,1,31,2,4,32,0,6,32,1,4,42,0,1,42,2,2,38,1,2,38,2,10,39,0,5,
/* out0330_em-eta10-phi16*/	8,31,0,2,31,1,1,31,2,12,103,0,1,103,2,1,27,1,1,38,0,7,38,2,6,
/* out0331_em-eta11-phi16*/	10,21,1,7,21,2,1,31,0,5,94,0,3,94,1,8,103,0,5,103,1,9,103,2,12,27,1,10,27,2,1,
/* out0332_em-eta12-phi16*/	7,21,0,4,21,1,5,21,2,1,94,0,11,94,2,1,27,0,8,27,1,1,
/* out0333_em-eta13-phi16*/	11,12,1,1,20,2,2,21,0,6,85,0,1,93,1,4,93,2,3,94,0,1,94,2,1,16,1,2,26,2,4,27,0,2,
/* out0334_em-eta14-phi16*/	7,12,1,3,20,2,4,85,0,2,93,2,6,16,1,3,26,0,1,26,2,3,
/* out0335_em-eta15-phi16*/	9,11,2,3,12,0,1,12,1,1,20,0,1,20,2,1,84,1,7,15,1,2,15,2,3,16,0,1,
/* out0336_em-eta16-phi16*/	6,11,2,6,84,0,2,84,1,2,84,2,2,15,1,1,15,2,3,
/* out0337_em-eta17-phi16*/	5,11,0,2,11,1,3,84,0,2,84,2,3,15,0,3,
/* out0338_em-eta18-phi16*/	2,11,1,1,15,0,3,
/* out0339_em-eta19-phi16*/	0,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	0,
/* out0343_em-eta3-phi17*/	0,
/* out0344_em-eta4-phi17*/	0,
/* out0345_em-eta5-phi17*/	8,52,1,6,52,2,9,53,0,12,53,1,8,53,2,4,64,0,1,64,1,2,64,2,4,
/* out0346_em-eta6-phi17*/	8,44,0,6,44,1,1,44,2,7,40,1,6,51,2,1,52,0,13,52,1,2,52,2,7,
/* out0347_em-eta7-phi17*/	12,33,0,1,33,1,15,43,2,5,44,0,6,44,1,12,44,2,8,39,1,1,39,2,1,40,0,7,40,1,10,51,0,1,51,2,4,
/* out0348_em-eta8-phi17*/	8,32,1,3,32,2,10,33,0,7,33,1,1,39,0,2,39,1,2,39,2,14,40,0,1,
/* out0349_em-eta9-phi17*/	6,22,1,3,32,0,10,32,2,6,28,1,9,39,0,7,39,2,1,
/* out0350_em-eta10-phi17*/	4,22,0,1,22,1,13,28,0,6,28,1,7,
/* out0351_em-eta11-phi17*/	9,21,2,5,22,0,7,94,1,8,94,2,1,95,0,12,95,1,8,95,2,4,27,2,10,28,0,2,
/* out0352_em-eta12-phi17*/	5,21,0,1,21,2,9,94,2,12,27,0,4,27,2,5,
/* out0353_em-eta13-phi17*/	7,12,1,5,21,0,4,85,0,2,85,1,8,94,2,1,16,1,7,27,0,1,
/* out0354_em-eta14-phi17*/	5,12,0,1,12,1,6,85,0,8,16,0,3,16,1,4,
/* out0355_em-eta15-phi17*/	6,12,0,5,84,1,4,84,2,1,85,0,3,15,2,2,16,0,4,
/* out0356_em-eta16-phi17*/	5,11,0,3,11,2,3,12,0,1,84,2,6,15,2,5,
/* out0357_em-eta17-phi17*/	4,11,0,10,84,2,4,15,0,1,15,2,3,
/* out0358_em-eta18-phi17*/	3,11,0,1,11,1,1,15,0,1,
/* out0359_em-eta19-phi17*/	0,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	0,
/* out0363_em-eta3-phi18*/	0,
/* out0364_em-eta4-phi18*/	0,
/* out0365_em-eta5-phi18*/	8,41,1,9,41,2,6,42,0,4,42,1,2,42,2,1,53,0,4,53,1,8,53,2,12,
/* out0366_em-eta6-phi18*/	8,34,0,7,34,1,1,34,2,6,30,1,1,40,2,6,41,0,13,41,1,7,41,2,2,
/* out0367_em-eta7-phi18*/	12,24,1,5,33,0,1,33,2,15,34,0,8,34,1,12,34,2,6,29,1,1,29,2,1,30,0,1,30,1,4,40,0,7,40,2,10,
/* out0368_em-eta8-phi18*/	8,23,1,10,23,2,3,33,0,7,33,2,1,29,0,2,29,1,14,29,2,2,40,0,1,
/* out0369_em-eta9-phi18*/	6,22,2,3,23,0,10,23,1,6,28,2,9,29,0,7,29,1,1,
/* out0370_em-eta10-phi18*/	4,22,0,1,22,2,13,28,0,6,28,2,7,
/* out0371_em-eta11-phi18*/	9,13,1,5,22,0,7,86,0,1,86,1,8,95,0,4,95,1,8,95,2,12,17,1,10,28,0,2,
/* out0372_em-eta12-phi18*/	5,13,0,1,13,1,9,86,0,12,17,0,4,17,1,5,
/* out0373_em-eta13-phi18*/	7,12,2,5,13,0,4,85,1,8,85,2,2,86,0,1,16,2,7,17,0,1,
/* out0374_em-eta14-phi18*/	5,12,0,1,12,2,6,85,2,8,16,0,3,16,2,4,
/* out0375_em-eta15-phi18*/	6,12,0,5,80,0,1,80,1,4,85,2,3,7,1,2,16,0,4,
/* out0376_em-eta16-phi18*/	5,5,1,1,5,2,3,12,0,1,80,0,6,7,1,5,
/* out0377_em-eta17-phi18*/	4,5,1,4,80,0,4,7,0,1,7,1,3,
/* out0378_em-eta18-phi18*/	2,5,1,2,7,0,1,
/* out0379_em-eta19-phi18*/	0,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	0,
/* out0383_em-eta3-phi19*/	0,
/* out0384_em-eta4-phi19*/	0,
/* out0385_em-eta5-phi19*/	6,31,1,12,31,2,1,41,2,4,42,0,12,42,1,14,42,2,15,
/* out0386_em-eta6-phi19*/	11,24,1,1,24,2,1,34,0,1,34,1,2,34,2,3,30,1,5,30,2,7,31,0,6,31,1,4,41,0,3,41,2,4,
/* out0387_em-eta7-phi19*/	9,24,0,5,24,1,10,24,2,10,34,1,1,34,2,1,29,2,1,30,0,13,30,1,6,30,2,4,
/* out0388_em-eta8-phi19*/	6,15,1,4,23,2,9,24,0,9,19,1,6,29,0,2,29,2,12,
/* out0389_em-eta9-phi19*/	9,14,1,4,14,2,1,15,0,1,15,1,2,23,0,6,23,2,4,18,1,10,18,2,2,29,0,5,
/* out0390_em-eta10-phi19*/	8,14,0,2,14,1,12,14,2,1,87,0,1,87,2,1,17,2,1,18,0,7,18,1,6,
/* out0391_em-eta11-phi19*/	10,13,1,1,13,2,7,14,0,5,86,1,8,86,2,3,87,0,12,87,1,9,87,2,5,17,1,1,17,2,10,
/* out0392_em-eta12-phi19*/	7,13,0,4,13,1,1,13,2,5,86,0,1,86,2,11,17,0,8,17,2,1,
/* out0393_em-eta13-phi19*/	11,6,1,2,12,2,1,13,0,6,81,0,3,81,1,4,85,2,1,86,0,1,86,2,1,8,1,4,16,2,2,17,0,2,
/* out0394_em-eta14-phi19*/	7,6,1,4,12,2,3,81,0,6,85,2,2,8,0,1,8,1,3,16,2,3,
/* out0395_em-eta15-phi19*/	9,5,2,3,6,0,1,6,1,1,12,0,1,12,2,1,80,1,7,7,1,3,7,2,2,16,0,1,
/* out0396_em-eta16-phi19*/	6,5,2,5,80,0,2,80,1,2,80,2,2,7,1,3,7,2,1,
/* out0397_em-eta17-phi19*/	4,5,1,4,80,0,3,80,2,2,7,0,3,
/* out0398_em-eta18-phi19*/	2,5,1,1,7,0,3,
/* out0399_em-eta19-phi19*/	0,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	0,
/* out0403_em-eta3-phi20*/	0,
/* out0404_em-eta4-phi20*/	0,
/* out0405_em-eta5-phi20*/	3,21,0,11,21,1,2,31,2,13,
/* out0406_em-eta6-phi20*/	7,20,1,11,20,2,3,21,0,2,21,2,1,30,2,2,31,0,10,31,2,2,
/* out0407_em-eta7-phi20*/	11,16,0,16,16,1,5,16,2,6,24,0,1,24,2,5,19,1,3,19,2,5,20,0,6,20,1,5,30,0,2,30,2,3,
/* out0408_em-eta8-phi20*/	8,15,0,1,15,1,9,15,2,10,16,2,1,24,0,1,19,0,8,19,1,7,19,2,5,
/* out0409_em-eta9-phi20*/	7,8,1,1,14,2,5,15,0,11,15,1,1,10,1,2,18,2,10,19,0,5,
/* out0410_em-eta10-phi20*/	10,8,1,1,14,0,5,14,2,9,82,1,1,87,0,2,87,1,2,87,2,4,9,1,2,18,0,8,18,2,4,
/* out0411_em-eta11-phi20*/	11,7,1,7,13,2,1,14,0,4,82,0,5,82,1,8,87,0,1,87,1,5,87,2,6,9,1,8,17,2,2,18,0,1,
/* out0412_em-eta12-phi20*/	13,7,0,2,7,1,5,13,0,1,13,2,3,81,1,3,82,0,8,86,2,1,8,1,2,8,2,2,9,0,2,9,1,2,17,0,1,17,2,2,
/* out0413_em-eta13-phi20*/	7,6,1,5,6,2,4,81,0,1,81,1,8,81,2,2,8,1,5,8,2,2,
/* out0414_em-eta14-phi20*/	7,6,0,2,6,1,4,6,2,1,81,0,5,81,2,4,8,0,5,8,1,2,
/* out0415_em-eta15-phi20*/	8,5,2,1,6,0,5,77,0,1,80,1,3,80,2,2,81,0,1,7,2,4,8,0,2,
/* out0416_em-eta16-phi20*/	4,5,0,4,5,2,4,80,2,6,7,2,5,
/* out0417_em-eta17-phi20*/	5,5,0,3,5,1,2,76,1,2,80,2,3,7,0,3,
/* out0418_em-eta18-phi20*/	4,5,1,1,76,1,3,0,1,1,7,0,3,
/* out0419_em-eta19-phi20*/	1,0,1,1,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	0,
/* out0423_em-eta3-phi21*/	0,
/* out0424_em-eta4-phi21*/	0,
/* out0425_em-eta5-phi21*/	4,13,0,2,21,0,3,21,1,14,21,2,7,
/* out0426_em-eta6-phi21*/	5,10,0,3,16,1,2,12,1,9,20,2,12,21,2,8,
/* out0427_em-eta7-phi21*/	10,9,1,3,9,2,1,10,0,5,16,1,9,16,2,8,11,1,10,11,2,1,19,2,1,20,0,10,20,2,1,
/* out0428_em-eta8-phi21*/	10,9,0,2,9,1,12,15,2,6,16,2,1,10,1,1,10,2,2,11,0,3,11,1,5,19,0,3,19,2,5,
/* out0429_em-eta9-phi21*/	7,8,1,8,8,2,5,9,0,1,15,0,3,10,0,2,10,1,11,10,2,3,
/* out0430_em-eta10-phi21*/	8,7,2,1,8,0,8,8,1,6,82,1,1,9,1,1,9,2,5,10,0,6,10,1,2,
/* out0431_em-eta11-phi21*/	8,7,1,3,7,2,9,79,0,1,82,1,6,82,2,8,9,0,3,9,1,3,9,2,5,
/* out0432_em-eta12-phi21*/	7,7,0,9,7,1,1,78,1,3,82,0,3,82,2,7,8,2,2,9,0,7,
/* out0433_em-eta13-phi21*/	7,1,1,1,6,2,6,7,0,2,78,0,4,81,1,1,81,2,5,8,2,8,
/* out0434_em-eta14-phi21*/	7,6,0,3,6,2,4,77,1,3,78,0,1,81,2,5,8,0,6,8,2,1,
/* out0435_em-eta15-phi21*/	7,0,1,2,6,0,4,77,0,3,77,1,4,1,1,3,7,2,1,8,0,1,
/* out0436_em-eta16-phi21*/	6,0,1,3,5,0,4,77,0,6,80,2,1,1,1,2,7,2,2,
/* out0437_em-eta17-phi21*/	12,0,0,1,0,1,1,5,0,5,5,1,1,76,1,3,76,2,3,0,1,1,0,2,1,1,0,1,1,1,1,7,0,2,7,2,1,
/* out0438_em-eta18-phi21*/	2,76,1,4,0,1,4,
/* out0439_em-eta19-phi21*/	1,0,1,2,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	0,
/* out0443_em-eta3-phi22*/	0,
/* out0444_em-eta4-phi22*/	0,
/* out0445_em-eta5-phi22*/	5,6,1,1,12,1,1,12,2,3,13,0,14,13,2,14,
/* out0446_em-eta6-phi22*/	5,10,0,2,6,1,1,12,0,10,12,1,6,12,2,12,
/* out0447_em-eta7-phi22*/	8,4,1,4,9,2,7,10,0,6,10,2,15,5,1,4,11,1,1,11,2,15,12,0,5,
/* out0448_em-eta8-phi22*/	8,3,1,1,4,1,1,9,0,10,9,1,1,9,2,8,4,1,5,10,2,2,11,0,13,
/* out0449_em-eta9-phi22*/	8,3,1,7,8,2,9,9,0,3,3,2,1,4,0,1,4,1,4,10,0,4,10,2,9,
/* out0450_em-eta10-phi22*/	8,2,1,5,2,2,1,3,0,3,8,0,8,8,2,2,3,1,8,9,2,1,10,0,4,
/* out0451_em-eta11-phi22*/	11,2,0,3,2,1,8,7,2,5,79,0,12,79,2,4,82,2,1,2,2,1,3,0,1,3,1,4,9,0,2,9,2,5,
/* out0452_em-eta12-phi22*/	10,1,1,4,1,2,4,2,0,1,7,0,3,7,2,1,78,1,10,79,2,2,2,1,7,2,2,1,9,0,2,
/* out0453_em-eta13-phi22*/	8,1,0,1,1,1,8,78,0,7,78,1,1,78,2,2,2,0,1,2,1,7,8,2,1,
/* out0454_em-eta14-phi22*/	12,0,1,1,0,2,2,1,0,3,1,1,2,6,0,1,6,2,1,77,1,5,78,0,3,1,1,2,1,2,3,2,0,4,8,0,1,
/* out0455_em-eta15-phi22*/	8,0,1,4,0,2,2,77,0,1,77,1,3,77,2,3,1,0,1,1,1,5,1,2,1,
/* out0456_em-eta16-phi22*/	7,0,0,1,0,1,4,0,2,1,77,0,4,77,2,2,1,0,2,1,1,3,
/* out0457_em-eta17-phi22*/	6,0,0,4,0,1,1,76,2,5,77,0,1,0,2,3,1,0,3,
/* out0458_em-eta18-phi22*/	4,76,1,3,76,2,3,0,1,2,0,2,3,
/* out0459_em-eta19-phi22*/	2,0,1,3,0,2,1,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	0,
/* out0463_em-eta3-phi23*/	0,
/* out0464_em-eta4-phi23*/	0,
/* out0465_em-eta5-phi23*/	4,6,0,4,6,1,8,6,2,16,13,2,2,
/* out0466_em-eta6-phi23*/	6,5,1,3,5,2,11,6,0,12,6,1,6,12,0,1,12,2,1,
/* out0467_em-eta7-phi23*/	7,4,0,7,4,1,9,4,2,16,10,2,1,5,0,14,5,1,9,5,2,5,
/* out0468_em-eta8-phi23*/	8,3,1,2,3,2,12,4,0,9,4,1,2,4,0,1,4,1,5,4,2,16,5,0,2,
/* out0469_em-eta9-phi23*/	6,3,0,9,3,1,6,3,2,4,3,2,6,4,0,14,4,1,2,
/* out0470_em-eta10-phi23*/	6,2,1,1,2,2,13,3,0,4,3,0,2,3,1,3,3,2,9,
/* out0471_em-eta11-phi23*/	8,2,0,9,2,1,2,2,2,2,79,0,3,79,2,9,2,2,2,3,0,13,3,1,1,
/* out0472_em-eta12-phi23*/	7,1,2,8,2,0,3,78,1,2,78,2,5,79,2,1,2,1,1,2,2,9,
/* out0473_em-eta13-phi23*/	7,1,0,6,1,1,1,1,2,4,78,2,8,2,0,8,2,1,1,2,2,3,
/* out0474_em-eta14-phi23*/	8,0,2,2,1,0,6,77,1,1,77,2,1,78,0,1,78,2,1,1,2,7,2,0,3,
/* out0475_em-eta15-phi23*/	4,0,2,7,77,2,6,1,0,1,1,2,5,
/* out0476_em-eta16-phi23*/	4,0,0,4,0,2,2,77,2,4,1,0,5,
/* out0477_em-eta17-phi23*/	4,0,0,5,76,2,1,0,2,2,1,0,3,
/* out0478_em-eta18-phi23*/	4,0,0,1,76,1,1,76,2,4,0,2,5,
/* out0479_em-eta19-phi23*/	2,0,1,2,0,2,1
};