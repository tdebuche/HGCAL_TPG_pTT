parameter integer matrixH [0:11645] = {
/* num inputs = 284(in0-in283) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 22 */
//* total number of input in adders 3721 */

/* out0000_em-eta0-phi0*/	0,
/* out0001_em-eta1-phi0*/	0,
/* out0002_em-eta2-phi0*/	2,151,0,7,151,1,6,
/* out0003_em-eta3-phi0*/	6,138,1,16,138,2,13,139,0,5,139,1,4,151,0,9,151,2,5,
/* out0004_em-eta4-phi0*/	7,125,1,16,125,2,11,126,0,2,126,1,2,138,2,3,139,0,11,139,2,2,
/* out0005_em-eta5-phi0*/	5,111,1,16,111,2,1,125,2,5,126,0,12,126,2,1,
/* out0006_em-eta6-phi0*/	3,98,1,8,111,2,15,112,0,10,
/* out0007_em-eta7-phi0*/	4,98,1,8,98,2,13,99,0,3,112,0,2,
/* out0008_em-eta8-phi0*/	6,85,1,10,98,2,3,99,0,5,214,0,9,214,1,1,273,2,3,
/* out0009_em-eta9-phi0*/	12,85,1,3,85,2,11,86,0,2,214,0,7,214,1,6,214,2,6,265,0,1,265,1,2,273,1,4,273,2,10,101,1,3,101,2,13,
/* out0010_em-eta10-phi0*/	11,67,1,12,85,2,1,86,0,2,205,0,8,205,1,1,214,2,7,265,0,12,265,1,1,93,0,8,93,1,3,101,1,1,
/* out0011_em-eta11-phi0*/	11,67,1,2,67,2,9,205,0,4,205,1,3,205,2,6,257,0,1,257,1,2,265,0,3,265,2,2,93,0,8,93,2,2,
/* out0012_em-eta12-phi0*/	10,48,4,15,49,0,3,49,1,4,67,2,3,68,0,4,196,0,6,205,2,6,257,0,9,85,0,7,85,1,1,
/* out0013_em-eta13-phi0*/	12,48,5,8,49,0,13,49,1,12,49,4,10,49,5,2,196,0,6,196,1,1,196,2,3,249,1,1,257,0,4,257,2,1,85,0,7,
/* out0014_em-eta14-phi0*/	9,49,2,10,49,3,4,49,4,6,49,5,4,187,0,1,196,2,8,249,0,5,77,0,2,77,1,1,
/* out0015_em-eta15-phi0*/	8,29,4,12,30,1,4,49,2,4,49,3,12,187,0,7,196,2,2,249,0,5,77,0,6,
/* out0016_em-eta16-phi0*/	8,29,5,3,30,0,12,30,1,12,30,4,1,187,0,3,187,2,3,249,0,1,77,0,3,
/* out0017_em-eta17-phi0*/	7,30,2,1,30,3,1,30,4,11,30,5,2,187,2,5,242,2,3,70,2,2,
/* out0018_em-eta18-phi0*/	8,13,3,2,30,2,8,30,3,4,187,2,2,242,0,1,242,2,1,70,0,1,70,2,3,
/* out0019_em-eta19-phi0*/	5,12,2,16,12,3,4,13,3,12,13,4,16,30,3,11,
/* out0020_em-eta0-phi1*/	0,
/* out0021_em-eta1-phi1*/	0,
/* out0022_em-eta2-phi1*/	4,151,1,10,152,1,1,161,1,8,161,2,14,
/* out0023_em-eta3-phi1*/	5,139,1,11,151,2,11,152,0,16,152,1,5,152,2,4,
/* out0024_em-eta4-phi1*/	5,126,1,8,139,1,1,139,2,14,140,0,13,140,1,2,
/* out0025_em-eta5-phi1*/	6,112,1,2,126,0,2,126,1,6,126,2,15,127,0,6,140,0,1,
/* out0026_em-eta6-phi1*/	4,112,0,4,112,1,13,112,2,8,127,0,1,
/* out0027_em-eta7-phi1*/	4,99,0,2,99,1,12,112,2,7,113,0,1,
/* out0028_em-eta8-phi1*/	10,85,1,2,99,0,6,99,1,1,99,2,10,214,1,1,222,1,1,222,2,9,273,1,1,273,2,2,274,0,1,
/* out0029_em-eta9-phi1*/	16,85,1,1,85,2,4,86,0,5,86,1,8,99,2,1,214,1,7,215,0,6,222,1,3,222,2,4,265,1,4,273,1,11,273,2,1,274,0,7,101,1,11,101,2,3,102,0,5,
/* out0030_em-eta10-phi1*/	15,67,1,1,86,0,7,86,2,5,205,0,4,205,1,3,214,1,1,214,2,3,215,0,4,215,2,7,265,1,9,265,2,7,93,1,13,93,2,1,101,1,1,102,0,3,
/* out0031_em-eta11-phi1*/	17,67,1,1,67,2,4,68,0,2,68,1,14,68,2,3,69,0,2,69,1,12,205,1,8,205,2,3,206,0,3,215,2,1,257,1,6,265,2,6,266,0,1,85,1,1,93,2,12,94,0,1,
/* out0032_em-eta12-phi1*/	17,48,4,1,68,0,10,68,1,2,68,2,11,68,3,10,69,3,1,196,0,2,196,1,2,205,1,1,205,2,1,206,0,2,206,2,3,257,0,2,257,1,6,257,2,3,85,0,1,85,1,11,
/* out0033_em-eta13-phi1*/	12,48,5,8,49,5,6,50,1,3,51,1,3,68,3,6,69,3,4,196,0,2,196,1,9,249,1,2,257,2,7,85,0,1,85,2,9,
/* out0034_em-eta14-phi1*/	12,49,2,2,49,5,4,50,0,6,50,1,11,187,0,1,196,1,3,196,2,3,197,0,1,249,0,2,249,1,6,77,1,6,85,2,2,
/* out0035_em-eta15-phi1*/	11,29,4,4,50,0,10,50,2,1,50,3,5,187,0,3,187,1,4,249,0,3,249,2,3,77,0,4,77,1,2,77,2,2,
/* out0036_em-eta16-phi1*/	12,29,5,12,30,0,4,30,4,1,30,5,2,50,3,2,187,0,1,187,1,5,187,2,1,242,2,3,249,2,3,77,0,1,77,2,4,
/* out0037_em-eta17-phi1*/	8,30,2,1,30,4,3,30,5,11,31,1,1,187,1,1,187,2,3,242,2,6,70,2,6,
/* out0038_em-eta18-phi1*/	8,12,3,1,13,3,1,30,2,6,31,0,6,187,2,1,242,0,2,70,0,3,70,2,2,
/* out0039_em-eta19-phi1*/	4,12,0,1,12,3,11,13,3,1,31,0,3,
/* out0040_em-eta0-phi2*/	0,
/* out0041_em-eta1-phi2*/	0,
/* out0042_em-eta2-phi2*/	6,152,1,1,161,1,8,161,2,2,162,0,7,162,1,16,162,2,5,
/* out0043_em-eta3-phi2*/	6,140,1,2,152,1,9,152,2,12,153,0,12,153,1,4,162,0,8,
/* out0044_em-eta4-phi2*/	6,140,0,2,140,1,12,140,2,14,141,0,5,153,0,4,153,2,1,
/* out0045_em-eta5-phi2*/	5,127,0,6,127,1,15,127,2,6,140,2,2,141,0,2,
/* out0046_em-eta6-phi2*/	6,112,1,1,112,2,1,113,0,4,113,1,9,127,0,3,127,2,8,
/* out0047_em-eta7-phi2*/	5,99,1,3,100,1,1,113,0,11,113,1,1,113,2,6,
/* out0048_em-eta8-phi2*/	9,99,2,5,100,0,9,100,1,2,222,1,7,222,2,3,223,0,8,274,1,7,280,0,1,280,1,1,
/* out0049_em-eta9-phi2*/	16,86,1,8,86,2,2,100,0,5,215,0,5,215,1,6,222,1,5,223,0,4,223,2,3,274,0,7,274,1,6,274,2,6,102,0,4,102,1,13,102,2,2,108,0,1,108,1,1,
/* out0050_em-eta10-phi2*/	15,68,4,2,86,2,9,87,0,3,215,0,1,215,1,8,215,2,6,265,2,1,266,0,3,266,1,6,274,0,1,274,2,4,93,2,1,94,1,3,102,0,4,102,2,9,
/* out0051_em-eta11-phi2*/	14,68,4,14,68,5,9,69,0,11,69,1,4,87,0,1,206,0,9,206,1,2,215,2,2,266,0,11,266,1,1,266,2,2,94,0,10,94,1,4,94,2,1,
/* out0052_em-eta12-phi2*/	20,68,2,2,69,0,3,69,2,4,69,3,4,69,4,16,69,5,5,206,0,2,206,1,2,206,2,7,257,1,2,257,2,3,258,0,2,258,1,1,266,0,1,266,2,1,85,1,3,85,2,1,86,1,1,94,0,5,94,2,2,
/* out0053_em-eta13-phi2*/	12,50,4,6,51,1,10,69,2,5,69,3,7,196,1,1,197,0,5,206,2,4,249,1,1,257,2,2,258,0,7,85,2,4,86,0,6,
/* out0054_em-eta14-phi2*/	12,50,1,2,50,2,8,51,0,10,51,1,3,51,4,1,197,0,6,197,2,2,249,1,6,249,2,1,258,0,1,77,1,5,86,0,4,
/* out0055_em-eta15-phi2*/	9,50,2,7,50,3,5,51,3,3,51,4,5,187,1,1,197,2,5,249,2,6,77,1,2,77,2,4,
/* out0056_em-eta16-phi2*/	15,29,5,1,30,5,1,31,1,1,32,1,4,50,3,4,51,3,8,187,1,3,188,1,1,242,0,1,242,2,2,249,2,2,250,0,1,70,2,1,77,2,5,78,0,1,
/* out0057_em-eta17-phi2*/	9,31,1,10,31,2,1,32,1,3,187,1,2,188,1,2,242,0,5,242,2,1,70,0,4,70,2,2,
/* out0058_em-eta18-phi2*/	8,31,0,4,31,1,4,31,2,3,31,3,1,187,2,1,188,1,1,242,0,1,70,0,3,
/* out0059_em-eta19-phi2*/	3,12,0,15,31,0,3,31,3,12,
/* out0060_em-eta0-phi3*/	0,
/* out0061_em-eta1-phi3*/	0,
/* out0062_em-eta2-phi3*/	4,162,2,10,163,0,6,163,1,11,170,0,3,
/* out0063_em-eta3-phi3*/	8,153,1,12,153,2,9,154,0,5,154,1,2,162,0,1,162,2,1,163,0,10,163,2,6,
/* out0064_em-eta4-phi3*/	5,141,0,5,141,1,16,141,2,5,153,2,6,154,0,6,
/* out0065_em-eta5-phi3*/	6,127,1,1,127,2,2,128,0,4,128,1,10,141,0,4,141,2,10,
/* out0066_em-eta6-phi3*/	5,113,1,6,113,2,1,114,1,1,128,0,12,128,2,5,
/* out0067_em-eta7-phi3*/	3,100,1,2,113,2,9,114,0,9,
/* out0068_em-eta8-phi3*/	10,100,0,1,100,1,10,100,2,6,114,0,1,223,0,2,223,1,7,274,1,1,280,0,12,280,1,7,280,2,9,
/* out0069_em-eta9-phi3*/	21,87,1,6,100,0,1,100,2,8,216,0,2,223,0,2,223,1,4,223,2,12,274,1,2,274,2,5,275,0,6,275,1,4,280,0,2,280,1,7,280,2,5,102,1,3,102,2,2,103,0,2,103,1,4,108,0,14,108,1,14,108,2,14,
/* out0070_em-eta10-phi3*/	12,87,0,8,87,1,3,87,2,1,215,1,2,216,0,12,216,2,2,266,1,8,274,2,1,275,0,7,94,1,3,102,2,3,103,0,11,
/* out0071_em-eta11-phi3*/	14,68,5,7,69,5,2,70,1,1,71,1,4,87,0,4,87,2,3,206,1,5,216,2,7,266,1,1,266,2,11,267,0,1,94,1,6,94,2,7,103,0,1,
/* out0072_em-eta12-phi3*/	13,69,2,5,69,5,9,70,0,5,70,1,14,71,1,1,206,1,7,206,2,1,207,0,3,258,1,9,266,2,2,86,1,5,94,2,6,95,0,1,
/* out0073_em-eta13-phi3*/	15,50,4,10,50,5,3,69,2,2,70,0,11,70,3,3,197,0,3,197,1,3,206,2,1,207,2,1,258,0,4,258,1,2,258,2,4,86,0,3,86,1,6,86,2,2,
/* out0074_em-eta14-phi3*/	12,50,5,10,51,0,6,51,4,4,51,5,4,197,0,1,197,1,5,197,2,2,250,1,2,258,0,2,258,2,3,86,0,3,86,2,5,
/* out0075_em-eta15-phi3*/	11,51,2,6,51,3,3,51,4,6,51,5,4,197,2,6,249,2,1,250,0,5,250,1,1,77,2,1,78,0,3,78,1,2,
/* out0076_em-eta16-phi3*/	9,31,4,6,32,1,4,51,2,5,51,3,2,188,1,1,188,2,4,242,0,1,250,0,5,78,0,6,
/* out0077_em-eta17-phi3*/	8,31,2,1,32,0,7,32,1,5,188,1,4,242,0,5,250,0,1,70,0,3,78,0,2,
/* out0078_em-eta18-phi3*/	5,31,2,8,32,0,2,32,4,2,188,1,2,70,0,2,
/* out0079_em-eta19-phi3*/	4,31,2,3,31,3,3,32,3,11,32,4,2,
/* out0080_em-eta0-phi4*/	0,
/* out0081_em-eta1-phi4*/	0,
/* out0082_em-eta2-phi4*/	7,163,1,5,163,2,3,164,0,2,164,1,9,170,0,13,170,1,16,170,2,16,
/* out0083_em-eta3-phi4*/	9,154,0,1,154,1,14,154,2,4,155,0,2,155,1,1,163,2,7,164,0,14,164,1,1,164,2,3,
/* out0084_em-eta4-phi4*/	6,141,2,1,142,0,4,142,1,13,154,0,4,154,2,12,155,0,4,
/* out0085_em-eta5-phi4*/	6,128,1,6,128,2,2,129,0,1,129,1,3,142,0,12,142,2,8,
/* out0086_em-eta6-phi4*/	3,114,1,7,128,2,9,129,0,10,
/* out0087_em-eta7-phi4*/	3,114,0,5,114,1,7,114,2,10,
/* out0088_em-eta8-phi4*/	14,100,1,1,100,2,2,101,0,5,101,1,6,114,0,1,114,2,3,223,1,2,224,0,2,224,1,2,280,0,1,280,1,1,280,2,2,281,0,2,281,2,1,
/* out0089_em-eta9-phi4*/	22,87,1,3,101,0,11,216,0,1,216,1,1,223,1,3,223,2,1,224,0,14,224,1,1,224,2,6,275,0,1,275,1,12,275,2,4,281,0,6,281,1,5,281,2,1,103,1,10,108,0,1,108,1,1,108,2,2,109,0,8,109,1,5,109,2,3,
/* out0090_em-eta10-phi4*/	13,87,1,4,87,2,8,88,0,1,216,0,1,216,1,13,216,2,1,224,2,1,267,1,4,275,0,2,275,2,10,103,0,2,103,1,2,103,2,13,
/* out0091_em-eta11-phi4*/	13,70,4,12,71,1,7,87,2,4,88,0,1,207,0,5,207,1,1,216,1,2,216,2,6,267,0,9,267,1,4,95,0,5,95,1,8,103,2,2,
/* out0092_em-eta12-phi4*/	15,70,1,1,70,2,11,70,5,1,71,0,13,71,1,4,71,4,4,207,0,8,207,1,1,207,2,2,258,1,4,267,0,6,267,2,1,86,1,1,95,0,10,95,2,1,
/* out0093_em-eta13-phi4*/	11,70,2,5,70,3,11,71,3,7,71,4,4,197,1,1,207,2,8,258,2,7,259,0,2,86,1,3,86,2,4,87,0,1,
/* out0094_em-eta14-phi4*/	14,50,5,3,51,5,6,52,1,6,53,1,4,70,3,2,71,3,3,197,1,5,198,0,3,250,1,5,258,2,2,259,0,1,78,1,2,86,2,5,87,0,2,
/* out0095_em-eta15-phi4*/	13,51,2,4,51,5,2,52,0,8,52,1,6,188,2,2,197,1,2,197,2,1,198,0,2,198,2,1,250,0,1,250,1,4,250,2,1,78,1,7,
/* out0096_em-eta16-phi4*/	9,31,4,9,51,2,1,52,0,6,188,2,6,250,0,2,250,2,3,78,0,2,78,1,1,78,2,3,
/* out0097_em-eta17-phi4*/	10,31,4,1,31,5,7,32,0,5,188,0,2,188,1,2,188,2,1,250,0,1,250,2,2,78,0,2,78,2,3,
/* out0098_em-eta18-phi4*/	4,32,0,2,32,4,9,32,5,1,188,1,2,
/* out0099_em-eta19-phi4*/	3,32,2,2,32,3,5,32,4,3,
/* out0100_em-eta0-phi5*/	0,
/* out0101_em-eta1-phi5*/	0,
/* out0102_em-eta2-phi5*/	4,164,1,6,164,2,1,165,0,1,165,1,3,
/* out0103_em-eta3-phi5*/	7,155,0,1,155,1,15,155,2,2,164,2,12,165,0,15,165,1,2,165,2,9,
/* out0104_em-eta4-phi5*/	6,142,1,3,142,2,2,143,0,2,143,1,8,155,0,9,155,2,14,
/* out0105_em-eta5-phi5*/	4,129,1,10,129,2,1,142,2,6,143,0,14,
/* out0106_em-eta6-phi5*/	4,115,1,2,129,0,5,129,1,3,129,2,15,
/* out0107_em-eta7-phi5*/	4,114,1,1,114,2,3,115,0,12,115,1,6,
/* out0108_em-eta8-phi5*/	4,101,1,10,101,2,4,115,0,4,224,1,3,
/* out0109_em-eta9-phi5*/	15,88,1,2,101,2,12,217,0,1,224,1,10,224,2,7,275,2,1,276,0,4,276,1,8,281,0,8,281,1,11,281,2,14,104,1,6,109,0,8,109,1,11,109,2,13,
/* out0110_em-eta10-phi5*/	10,88,0,6,88,1,6,217,0,13,224,2,2,267,1,3,275,2,1,276,0,12,103,2,1,104,0,13,104,1,2,
/* out0111_em-eta11-phi5*/	11,70,4,4,70,5,6,88,0,8,207,1,3,217,0,2,217,2,8,267,1,5,267,2,9,95,1,8,95,2,4,104,0,3,
/* out0112_em-eta12-phi5*/	10,70,5,9,71,0,3,71,2,1,71,4,6,71,5,15,207,1,10,259,1,5,267,2,6,87,1,1,95,2,11,
/* out0113_em-eta13-phi5*/	12,52,4,4,71,2,15,71,3,6,71,4,2,71,5,1,198,0,3,207,1,1,207,2,5,259,0,7,259,1,3,87,0,3,87,1,7,
/* out0114_em-eta14-phi5*/	9,52,1,1,52,2,1,52,4,4,53,0,6,53,1,12,198,0,7,250,1,2,259,0,6,87,0,8,
/* out0115_em-eta15-phi5*/	12,52,0,1,52,1,3,52,2,14,52,3,1,53,0,2,198,0,1,198,2,5,250,1,2,250,2,4,78,1,4,78,2,2,87,0,2,
/* out0116_em-eta16-phi5*/	9,31,5,1,52,0,1,52,2,1,52,3,13,188,0,1,188,2,3,198,2,2,250,2,5,78,2,6,
/* out0117_em-eta17-phi5*/	6,31,5,8,32,5,5,52,3,2,188,0,10,250,2,1,78,2,2,
/* out0118_em-eta18-phi5*/	5,32,2,2,32,5,10,33,0,1,188,0,3,188,1,1,
/* out0119_em-eta19-phi5*/	2,32,2,12,33,0,1,
/* out0120_em-eta0-phi6*/	0,
/* out0121_em-eta1-phi6*/	0,
/* out0122_em-eta2-phi6*/	3,165,1,3,166,0,1,166,1,6,
/* out0123_em-eta3-phi6*/	6,156,0,2,156,1,15,156,2,1,165,1,8,165,2,7,166,0,12,
/* out0124_em-eta4-phi6*/	6,143,1,8,143,2,2,144,0,2,144,1,3,156,0,14,156,2,9,
/* out0125_em-eta5-phi6*/	4,130,0,1,130,1,10,143,2,14,144,0,6,
/* out0126_em-eta6-phi6*/	4,115,1,2,130,0,15,130,1,3,130,2,5,
/* out0127_em-eta7-phi6*/	4,115,1,6,115,2,12,116,0,3,116,1,1,
/* out0128_em-eta8-phi6*/	5,102,0,4,102,1,10,115,2,4,225,0,1,225,1,3,
/* out0129_em-eta9-phi6*/	16,88,1,2,102,0,12,217,1,1,225,0,15,225,1,3,225,2,8,276,1,8,276,2,4,277,0,1,282,0,14,282,1,11,282,2,8,104,1,6,110,0,13,110,1,11,110,2,8,
/* out0130_em-eta10-phi6*/	10,88,1,6,88,2,6,217,1,13,225,2,2,268,1,3,276,2,12,277,0,1,104,1,2,104,2,13,105,0,1,
/* out0131_em-eta11-phi6*/	11,72,4,4,73,1,6,88,2,8,208,0,3,217,1,2,217,2,8,268,0,9,268,1,5,96,0,4,96,1,8,104,2,3,
/* out0132_em-eta12-phi6*/	10,72,0,1,72,1,15,72,2,6,73,0,3,73,1,9,208,0,10,259,1,5,268,0,6,87,1,1,96,0,11,
/* out0133_em-eta13-phi6*/	12,52,4,4,72,0,15,72,1,1,72,2,2,72,3,6,198,1,3,208,0,1,208,2,5,259,1,3,259,2,7,87,1,7,87,2,3,
/* out0134_em-eta14-phi6*/	9,52,4,4,52,5,12,53,0,6,53,4,1,53,5,1,198,1,7,251,1,2,259,2,6,87,2,8,
/* out0135_em-eta15-phi6*/	12,53,0,2,53,2,1,53,3,1,53,4,14,53,5,2,198,1,1,198,2,5,251,0,4,251,1,2,79,0,2,79,1,4,87,2,2,
/* out0136_em-eta16-phi6*/	9,34,1,1,53,2,1,53,3,13,53,4,1,189,1,1,189,2,3,198,2,2,251,0,5,79,0,6,
/* out0137_em-eta17-phi6*/	6,33,1,5,34,1,8,53,3,2,189,1,4,251,0,1,79,0,2,
/* out0138_em-eta18-phi6*/	3,33,0,2,33,1,10,189,1,2,
/* out0139_em-eta19-phi6*/	1,33,0,10,
/* out0140_em-eta0-phi7*/	0,
/* out0141_em-eta1-phi7*/	0,
/* out0142_em-eta2-phi7*/	7,166,1,9,166,2,2,167,0,3,167,1,5,171,0,16,171,1,15,171,2,16,
/* out0143_em-eta3-phi7*/	9,156,1,1,156,2,2,157,0,4,157,1,14,157,2,1,166,0,3,166,1,1,166,2,14,167,0,7,
/* out0144_em-eta4-phi7*/	6,144,1,13,144,2,4,145,0,1,156,2,4,157,0,12,157,2,4,
/* out0145_em-eta5-phi7*/	6,130,1,3,130,2,1,131,0,2,131,1,6,144,0,8,144,2,12,
/* out0146_em-eta6-phi7*/	3,116,1,7,130,2,10,131,0,9,
/* out0147_em-eta7-phi7*/	3,116,0,10,116,1,7,116,2,5,
/* out0148_em-eta8-phi7*/	14,102,1,6,102,2,5,103,0,2,103,1,1,116,0,3,116,2,1,225,1,3,226,0,3,226,1,1,282,0,1,282,2,2,283,0,2,283,1,1,283,2,1,
/* out0149_em-eta9-phi7*/	20,89,1,3,102,2,11,218,0,1,218,1,1,225,1,7,225,2,5,226,0,7,277,0,4,277,1,12,277,2,1,282,0,1,282,1,5,282,2,6,105,1,10,110,0,3,110,1,5,110,2,8,111,0,2,111,1,1,111,2,1,
/* out0150_em-eta10-phi7*/	13,88,2,1,89,0,8,89,1,4,218,0,13,218,1,1,218,2,1,225,2,1,268,1,4,277,0,10,277,2,1,105,0,13,105,1,2,105,2,2,
/* out0151_em-eta11-phi7*/	13,72,4,12,72,5,7,88,2,1,89,0,4,208,0,1,208,1,5,218,0,2,218,2,6,268,1,4,268,2,9,96,1,8,96,2,5,105,0,2,
/* out0152_em-eta12-phi7*/	15,72,2,4,72,5,4,73,0,13,73,1,1,73,4,11,73,5,1,208,0,1,208,1,8,208,2,2,260,1,4,268,0,1,268,2,6,88,1,1,96,0,1,96,2,10,
/* out0153_em-eta13-phi7*/	11,72,2,4,72,3,7,73,3,11,73,4,5,199,0,1,208,2,8,259,2,2,260,0,7,87,2,1,88,0,4,88,1,3,
/* out0154_em-eta14-phi7*/	14,52,5,4,53,5,7,54,1,6,55,1,3,72,3,3,73,3,2,198,1,3,199,0,5,251,1,5,259,2,1,260,0,2,79,1,2,87,2,2,88,0,5,
/* out0155_em-eta15-phi7*/	13,53,2,8,53,5,6,54,0,4,54,1,2,189,2,1,198,1,2,198,2,1,199,0,2,199,2,1,251,0,1,251,1,4,251,2,1,79,1,7,
/* out0156_em-eta16-phi7*/	9,33,4,9,53,2,6,54,0,1,189,2,6,251,0,3,251,2,2,79,0,3,79,1,1,79,2,2,
/* out0157_em-eta17-phi7*/	9,33,4,1,34,0,5,34,1,7,189,1,3,189,2,1,251,0,2,251,2,1,79,0,3,79,2,2,
/* out0158_em-eta18-phi7*/	4,33,1,1,33,2,9,34,0,2,189,1,2,
/* out0159_em-eta19-phi7*/	3,33,0,2,33,2,3,33,3,5,
/* out0160_em-eta0-phi8*/	0,
/* out0161_em-eta1-phi8*/	0,
/* out0162_em-eta2-phi8*/	4,167,1,11,167,2,6,168,1,10,171,1,1,
/* out0163_em-eta3-phi8*/	8,157,1,2,157,2,5,158,0,9,158,1,12,167,0,6,167,2,10,168,0,1,168,1,1,
/* out0164_em-eta4-phi8*/	5,145,0,5,145,1,16,145,2,5,157,2,6,158,0,6,
/* out0165_em-eta5-phi8*/	6,131,1,10,131,2,4,132,0,2,132,1,1,145,0,10,145,2,4,
/* out0166_em-eta6-phi8*/	5,116,1,1,117,0,1,117,1,6,131,0,5,131,2,12,
/* out0167_em-eta7-phi8*/	3,103,1,2,116,2,9,117,0,9,
/* out0168_em-eta8-phi8*/	9,103,0,6,103,1,10,103,2,1,116,2,1,226,1,8,278,1,1,283,0,9,283,1,7,283,2,12,
/* out0169_em-eta9-phi8*/	21,89,1,6,103,0,8,103,2,1,218,1,2,226,0,6,226,1,2,226,2,13,277,1,4,277,2,7,278,0,5,278,1,2,283,0,5,283,1,7,283,2,2,105,1,4,105,2,2,106,0,2,106,1,3,111,0,14,111,1,14,111,2,14,
/* out0170_em-eta10-phi8*/	12,89,0,1,89,1,3,89,2,8,218,1,12,218,2,2,219,0,2,269,1,8,277,2,7,278,0,1,97,1,3,105,2,11,106,0,3,
/* out0171_em-eta11-phi8*/	14,72,5,4,73,5,1,74,1,2,75,1,7,89,0,3,89,2,4,209,0,5,218,2,7,268,2,1,269,0,11,269,1,1,97,0,7,97,1,6,105,2,1,
/* out0172_em-eta12-phi8*/	13,72,5,1,73,2,5,73,5,14,74,0,5,74,1,9,208,1,3,209,0,7,209,2,1,260,1,9,269,0,2,88,1,5,96,2,1,97,0,6,
/* out0173_em-eta13-phi8*/	15,54,4,10,55,1,3,73,2,11,73,3,3,74,0,2,199,0,3,199,1,3,208,2,1,209,2,1,260,0,4,260,1,2,260,2,4,88,0,2,88,1,6,88,2,3,
/* out0174_em-eta14-phi8*/	12,54,1,4,54,2,4,55,0,6,55,1,10,199,0,5,199,1,1,199,2,2,251,1,2,260,0,3,260,2,2,88,0,5,88,2,3,
/* out0175_em-eta15-phi8*/	11,54,0,6,54,1,4,54,2,6,54,3,3,199,2,6,251,1,1,251,2,5,252,0,1,79,1,2,79,2,3,80,0,1,
/* out0176_em-eta16-phi8*/	9,33,4,6,33,5,4,54,0,5,54,3,2,189,0,2,189,2,5,243,1,1,251,2,5,79,2,6,
/* out0177_em-eta17-phi8*/	9,33,5,5,34,0,7,34,4,1,189,0,5,189,1,2,243,1,5,251,2,1,71,1,3,79,2,2,
/* out0178_em-eta18-phi8*/	5,33,2,2,34,0,2,34,4,8,189,1,1,71,1,2,
/* out0179_em-eta19-phi8*/	4,33,2,2,33,3,11,34,3,3,34,4,3,
/* out0180_em-eta0-phi9*/	0,
/* out0181_em-eta1-phi9*/	0,
/* out0182_em-eta2-phi9*/	6,159,1,1,168,0,7,168,1,5,168,2,16,169,0,9,169,2,1,
/* out0183_em-eta3-phi9*/	6,146,1,2,158,1,4,158,2,12,159,0,12,159,1,9,168,0,8,
/* out0184_em-eta4-phi9*/	6,145,2,5,146,0,14,146,1,12,146,2,2,158,0,1,158,2,4,
/* out0185_em-eta5-phi9*/	5,132,0,6,132,1,15,132,2,6,145,2,2,146,0,2,
/* out0186_em-eta6-phi9*/	6,117,1,9,117,2,4,118,0,1,118,1,1,132,0,8,132,2,3,
/* out0187_em-eta7-phi9*/	5,103,1,1,104,1,3,117,0,6,117,1,1,117,2,11,
/* out0188_em-eta8-phi9*/	9,103,1,2,103,2,9,104,0,5,104,1,1,226,1,3,227,0,10,278,1,7,283,1,1,283,2,1,
/* out0189_em-eta9-phi9*/	17,90,0,2,90,1,8,103,2,5,219,0,6,219,1,5,226,1,2,226,2,3,227,0,2,227,2,3,278,0,6,278,1,6,278,2,7,106,0,2,106,1,13,106,2,4,111,1,1,111,2,1,
/* out0190_em-eta10-phi9*/	15,74,4,2,89,2,3,90,0,9,219,0,8,219,1,1,219,2,6,269,1,6,269,2,3,270,0,1,278,0,4,278,2,1,97,1,3,98,0,1,106,0,9,106,2,4,
/* out0191_em-eta11-phi9*/	14,74,4,14,74,5,4,75,0,11,75,1,9,89,2,1,209,0,2,209,1,9,219,2,2,269,0,2,269,1,1,269,2,11,97,0,1,97,1,4,97,2,10,
/* out0192_em-eta12-phi9*/	20,74,0,4,74,1,5,74,2,16,74,3,4,75,0,3,75,4,2,209,0,2,209,1,2,209,2,7,260,1,1,260,2,2,261,0,3,261,1,2,269,0,1,269,2,1,88,1,1,89,0,1,89,1,3,97,0,2,97,2,5,
/* out0193_em-eta13-phi9*/	11,54,4,6,54,5,10,74,0,5,74,3,7,199,1,5,209,2,4,252,1,1,260,2,7,261,0,2,88,2,6,89,0,4,
/* out0194_em-eta14-phi9*/	12,54,2,1,54,5,3,55,0,10,55,4,8,55,5,2,199,1,6,199,2,2,252,0,1,252,1,6,260,2,1,80,1,5,88,2,4,
/* out0195_em-eta15-phi9*/	9,54,2,5,54,3,3,55,3,5,55,4,7,190,0,1,199,2,5,252,0,6,80,0,4,80,1,2,
/* out0196_em-eta16-phi9*/	15,33,5,4,34,5,1,35,1,1,36,1,1,54,3,8,55,3,4,189,0,3,190,0,3,243,1,1,243,2,2,251,2,1,252,0,2,71,2,1,79,2,1,80,0,5,
/* out0197_em-eta17-phi9*/	9,33,5,3,34,4,1,34,5,10,189,0,6,190,0,2,243,1,5,243,2,1,71,1,4,71,2,2,
/* out0198_em-eta18-phi9*/	7,34,2,4,34,3,1,34,4,3,34,5,4,189,1,1,243,1,1,71,1,3,
/* out0199_em-eta19-phi9*/	3,14,4,15,34,2,3,34,3,12,
/* out0200_em-eta0-phi10*/	0,
/* out0201_em-eta1-phi10*/	0,
/* out0202_em-eta2-phi10*/	4,159,1,1,160,1,10,169,0,7,169,2,15,
/* out0203_em-eta3-phi10*/	5,147,1,11,159,0,4,159,1,5,159,2,16,160,0,11,
/* out0204_em-eta4-phi10*/	5,133,1,8,146,1,2,146,2,13,147,0,14,147,1,1,
/* out0205_em-eta5-phi10*/	6,118,1,2,132,2,6,133,0,15,133,1,6,133,2,2,146,2,1,
/* out0206_em-eta6-phi10*/	4,118,0,8,118,1,13,118,2,4,132,2,1,
/* out0207_em-eta7-phi10*/	4,104,1,11,104,2,2,117,2,1,118,0,7,
/* out0208_em-eta8-phi10*/	8,104,0,10,104,1,1,104,2,6,220,0,1,227,0,4,227,2,6,278,2,1,279,0,4,
/* out0209_em-eta9-phi10*/	13,90,1,8,90,2,5,104,0,1,219,1,6,220,0,7,227,2,7,270,1,4,278,2,7,279,0,8,279,2,4,106,2,5,107,0,12,107,2,3,
/* out0210_em-eta10-phi10*/	13,76,1,1,90,0,5,90,2,7,210,0,3,219,1,4,219,2,7,220,0,1,270,0,7,270,1,9,98,0,1,98,1,13,106,2,3,107,2,1,
/* out0211_em-eta11-phi10*/	15,74,5,12,75,0,2,75,2,2,75,4,3,75,5,14,76,0,1,209,1,3,210,0,8,219,2,1,261,1,6,269,2,1,270,0,6,89,1,1,97,2,1,98,0,12,
/* out0212_em-eta12-phi10*/	17,56,4,1,74,3,1,75,2,10,75,3,10,75,4,11,75,5,2,200,0,2,200,1,1,209,1,2,209,2,3,210,0,1,210,2,1,261,0,3,261,1,6,261,2,2,89,1,11,89,2,1,
/* out0213_em-eta13-phi10*/	11,54,5,3,55,5,3,56,1,6,57,1,8,74,3,4,75,3,6,200,0,9,252,1,2,261,0,7,89,0,9,89,2,1,
/* out0214_em-eta14-phi10*/	11,55,2,6,55,5,11,56,0,2,56,1,4,199,1,1,200,0,4,200,2,2,252,1,6,252,2,2,80,1,6,89,0,2,
/* out0215_em-eta15-phi10*/	11,35,4,4,55,2,10,55,3,5,55,4,1,190,0,4,190,1,3,252,0,3,252,2,3,80,0,2,80,1,2,80,2,4,
/* out0216_em-eta16-phi10*/	8,35,1,2,36,1,12,55,3,2,190,0,5,243,2,3,252,0,3,80,0,4,80,2,1,
/* out0217_em-eta17-phi10*/	7,34,5,1,35,0,1,35,1,11,190,0,1,190,2,3,243,2,6,71,2,6,
/* out0218_em-eta18-phi10*/	7,14,5,1,34,2,6,35,0,6,190,2,1,243,1,2,71,1,3,71,2,2,
/* out0219_em-eta19-phi10*/	4,14,4,1,14,5,11,15,5,1,34,2,3,
/* out0220_em-eta0-phi11*/	0,
/* out0221_em-eta1-phi11*/	0,
/* out0222_em-eta2-phi11*/	2,160,1,6,160,2,7,
/* out0223_em-eta3-phi11*/	5,147,1,4,147,2,5,148,2,3,160,0,5,160,2,9,
/* out0224_em-eta4-phi11*/	7,133,1,2,133,2,2,134,0,7,134,1,12,147,0,2,147,2,11,148,2,2,
/* out0225_em-eta5-phi11*/	5,119,0,1,119,1,12,133,0,1,133,2,12,134,0,5,
/* out0226_em-eta6-phi11*/	3,105,1,4,118,2,10,119,0,11,
/* out0227_em-eta7-phi11*/	4,104,2,3,105,0,9,105,1,8,118,2,2,
/* out0228_em-eta8-phi11*/	6,91,1,10,104,2,5,105,0,3,220,0,1,220,1,5,279,0,2,
/* out0229_em-eta9-phi11*/	15,90,2,2,91,0,11,91,1,2,220,0,6,220,1,7,220,2,5,270,1,2,270,2,1,271,0,2,271,1,4,279,0,2,279,2,12,99,1,3,107,0,4,107,2,11,
/* out0230_em-eta10-phi11*/	15,76,1,9,90,2,2,91,0,1,210,0,1,210,1,8,220,2,7,262,1,1,270,1,1,270,2,12,271,0,2,98,1,3,98,2,8,99,0,4,99,1,1,107,2,1,
/* out0231_em-eta11-phi11*/	14,76,0,8,76,1,2,210,0,3,210,1,4,210,2,6,261,1,2,261,2,1,262,0,2,262,1,3,270,0,2,270,2,3,90,1,4,98,0,2,98,2,8,
/* out0232_em-eta12-phi11*/	11,56,4,15,56,5,4,75,2,4,76,0,3,200,1,5,210,2,5,261,2,9,262,0,2,89,1,1,89,2,7,90,0,4,
/* out0233_em-eta13-phi11*/	14,56,1,2,56,2,6,57,0,12,57,1,8,200,0,1,200,1,6,200,2,2,252,1,1,253,0,1,253,1,4,261,0,1,261,2,4,81,1,2,89,2,7,
/* out0234_em-eta14-phi11*/	11,56,0,10,56,1,4,56,2,6,56,3,4,200,2,8,252,2,5,253,0,3,80,1,1,80,2,2,81,0,3,81,1,2,
/* out0235_em-eta15-phi11*/	8,35,4,12,35,5,4,56,0,4,190,1,6,244,1,1,252,2,5,80,2,6,81,0,1,
/* out0236_em-eta16-phi11*/	10,35,2,1,36,0,12,36,1,3,190,1,3,190,2,3,244,0,1,244,1,3,252,2,1,72,1,3,80,2,3,
/* out0237_em-eta17-phi11*/	8,35,0,1,35,1,2,35,2,11,190,2,4,243,2,3,244,0,3,71,2,2,72,0,3,
/* out0238_em-eta18-phi11*/	8,35,0,8,35,3,4,190,2,1,243,1,1,243,2,1,71,1,1,71,2,3,72,0,1,
/* out0239_em-eta19-phi11*/	4,14,5,4,15,0,16,15,4,12,15,5,11,
/* out0240_em-eta0-phi12*/	0,
/* out0241_em-eta1-phi12*/	0,
/* out0242_em-eta2-phi12*/	1,149,1,13,
/* out0243_em-eta3-phi12*/	5,135,1,9,148,1,16,148,2,9,149,0,13,149,1,1,
/* out0244_em-eta4-phi12*/	7,120,1,4,134,0,1,134,1,4,134,2,14,135,0,10,135,1,3,148,2,2,
/* out0245_em-eta5-phi12*/	6,119,1,4,119,2,9,120,0,8,120,1,5,134,0,3,134,2,2,
/* out0246_em-eta6-phi12*/	6,105,1,3,105,2,1,106,0,4,106,1,6,119,0,4,119,2,7,
/* out0247_em-eta7-phi12*/	5,92,1,2,105,0,2,105,1,1,105,2,14,106,0,2,
/* out0248_em-eta8-phi12*/	8,91,1,4,91,2,6,92,0,3,92,1,2,105,0,2,105,2,1,221,0,8,271,1,2,
/* out0249_em-eta9-phi12*/	14,77,1,2,91,0,3,91,2,10,211,0,3,211,1,3,220,1,4,220,2,3,221,0,5,221,2,4,271,0,3,271,1,10,271,2,6,99,1,11,99,2,4,
/* out0250_em-eta10-phi12*/	14,76,1,4,76,2,5,77,0,2,91,0,1,210,1,1,211,0,12,211,2,1,220,2,1,262,1,6,271,0,9,271,2,1,99,0,12,99,1,1,99,2,4,
/* out0251_em-eta11-phi12*/	13,76,0,2,76,2,8,201,0,3,201,1,2,210,1,3,210,2,3,211,0,1,211,2,1,262,0,4,262,1,6,262,2,3,90,1,12,90,2,2,
/* out0252_em-eta12-phi12*/	13,56,5,12,57,5,7,58,1,2,59,1,2,76,0,2,76,2,1,200,1,1,201,0,9,210,2,1,253,1,3,262,0,7,90,0,10,90,2,1,
/* out0253_em-eta13-phi12*/	16,56,2,1,57,0,4,57,2,1,57,3,2,57,4,14,57,5,7,191,0,1,200,1,3,200,2,2,201,0,2,201,2,1,253,0,1,253,1,8,253,2,1,81,1,9,90,0,1,
/* out0254_em-eta14-phi12*/	10,56,2,3,56,3,8,57,3,10,57,4,2,191,0,5,200,2,2,253,0,8,81,0,6,81,1,2,81,2,1,
/* out0255_em-eta15-phi12*/	9,35,5,12,36,5,4,56,3,4,190,1,2,191,0,4,244,1,5,253,0,1,72,1,3,81,0,4,
/* out0256_em-eta16-phi12*/	10,36,0,4,36,4,9,36,5,3,181,1,1,190,1,2,190,2,2,191,0,1,244,0,1,244,1,4,72,1,6,
/* out0257_em-eta17-phi12*/	8,35,2,4,36,3,3,36,4,7,181,1,3,190,2,2,244,0,5,72,0,4,72,1,1,
/* out0258_em-eta18-phi12*/	5,35,3,11,36,3,1,181,1,1,244,0,2,72,0,4,
/* out0259_em-eta19-phi12*/	4,15,2,8,15,3,1,15,4,4,15,5,4,
/* out0260_em-eta0-phi13*/	0,
/* out0261_em-eta1-phi13*/	0,
/* out0262_em-eta2-phi13*/	5,136,1,1,149,1,2,149,2,8,150,0,14,150,2,8,
/* out0263_em-eta3-phi13*/	6,135,1,4,135,2,7,136,0,12,136,1,13,149,0,3,149,2,8,
/* out0264_em-eta4-phi13*/	6,120,1,5,120,2,3,121,0,6,121,1,9,135,0,6,135,2,9,
/* out0265_em-eta5-phi13*/	7,106,1,2,107,0,1,107,1,4,120,0,8,120,1,2,120,2,13,121,0,1,
/* out0266_em-eta6-phi13*/	4,106,0,4,106,1,8,106,2,13,107,0,1,
/* out0267_em-eta7-phi13*/	4,92,1,10,92,2,4,106,0,6,106,2,1,
/* out0268_em-eta8-phi13*/	7,92,0,12,92,1,2,92,2,4,212,0,2,221,0,3,221,2,5,272,0,5,
/* out0269_em-eta9-phi13*/	13,77,1,13,77,2,1,92,0,1,211,1,7,212,0,6,221,2,7,263,1,4,271,2,7,272,0,8,272,2,4,99,2,3,100,0,13,100,2,4,
/* out0270_em-eta10-phi13*/	10,77,0,11,211,1,6,211,2,9,262,2,1,263,0,5,263,1,7,271,2,2,91,0,1,91,1,10,99,2,5,
/* out0271_em-eta11-phi13*/	14,58,4,16,58,5,4,59,0,5,59,1,8,76,2,2,201,1,8,202,0,1,211,2,4,254,1,2,262,2,9,263,0,3,82,1,1,90,2,7,91,0,7,
/* out0272_em-eta12-phi13*/	18,57,5,1,58,0,2,58,1,14,58,2,7,59,0,4,59,1,6,201,0,2,201,1,3,201,2,5,253,1,1,253,2,1,254,0,2,254,1,4,262,0,1,262,2,3,82,1,5,90,0,1,90,2,6,
/* out0273_em-eta13-phi13*/	11,37,4,5,57,2,13,57,5,1,58,0,10,191,1,4,201,2,5,253,2,8,254,0,1,81,1,1,81,2,6,82,0,3,
/* out0274_em-eta14-phi13*/	10,37,4,5,38,1,13,57,2,2,57,3,4,191,0,2,191,1,5,245,1,1,253,0,2,253,2,5,81,2,8,
/* out0275_em-eta15-phi13*/	15,36,5,4,37,0,1,37,1,13,38,1,2,191,0,3,191,2,4,244,1,3,244,2,3,245,0,1,72,1,2,72,2,1,73,0,1,73,1,1,81,0,2,81,2,1,
/* out0276_em-eta16-phi13*/	9,36,2,10,36,5,5,37,0,2,181,1,1,181,2,3,191,2,2,244,2,5,72,1,1,72,2,4,
/* out0277_em-eta17-phi13*/	9,16,4,1,36,2,5,36,3,7,181,1,5,181,2,1,244,0,2,244,2,2,72,0,1,72,2,4,
/* out0278_em-eta18-phi13*/	6,17,1,5,35,3,1,36,3,5,181,1,1,244,0,2,72,0,3,
/* out0279_em-eta19-phi13*/	3,15,2,8,15,3,14,16,1,3,
/* out0280_em-eta0-phi14*/	0,
/* out0281_em-eta1-phi14*/	0,
/* out0282_em-eta2-phi14*/	7,136,1,1,136,2,1,137,0,7,137,1,16,137,2,5,150,0,2,150,2,8,
/* out0283_em-eta3-phi14*/	7,121,1,1,122,0,4,122,1,12,136,0,4,136,1,1,136,2,15,137,0,8,
/* out0284_em-eta4-phi14*/	5,108,1,5,121,0,7,121,1,6,121,2,16,122,0,5,
/* out0285_em-eta5-phi14*/	5,107,0,4,107,1,12,107,2,12,108,0,2,121,0,2,
/* out0286_em-eta6-phi14*/	5,93,1,12,93,2,1,106,2,2,107,0,10,107,2,1,
/* out0287_em-eta7-phi14*/	5,78,1,1,92,2,3,93,0,13,93,1,4,93,2,1,
/* out0288_em-eta8-phi14*/	10,78,0,2,78,1,10,92,2,5,212,0,1,212,1,10,213,0,1,213,1,1,264,0,4,272,0,3,272,2,4,
/* out0289_em-eta9-phi14*/	16,77,1,1,77,2,9,78,0,5,212,0,7,212,1,3,212,2,9,263,1,3,263,2,3,264,0,9,264,2,3,272,2,8,91,1,1,92,0,13,92,2,2,100,0,3,100,2,12,
/* out0290_em-eta10-phi14*/	16,58,5,1,59,5,1,60,1,3,77,0,3,77,2,6,202,0,6,202,1,7,211,2,1,212,2,2,263,0,4,263,1,2,263,2,10,91,0,1,91,1,5,91,2,11,92,2,1,
/* out0291_em-eta11-phi14*/	16,58,5,11,59,0,6,59,2,1,59,4,6,59,5,15,201,1,1,202,0,9,202,2,2,254,1,7,254,2,2,263,0,4,263,2,1,82,1,3,82,2,1,91,0,7,91,2,3,
/* out0292_em-eta12-phi14*/	16,58,2,9,58,3,6,59,0,1,59,3,7,59,4,10,192,0,4,192,1,1,201,1,2,201,2,4,202,2,1,254,0,5,254,1,3,254,2,2,82,0,1,82,1,7,82,2,3,
/* out0293_em-eta13-phi14*/	11,37,4,5,37,5,11,58,0,4,58,3,9,191,1,2,192,0,6,201,2,1,245,1,3,253,2,1,254,0,6,82,0,10,
/* out0294_em-eta14-phi14*/	10,37,2,1,37,4,1,37,5,3,38,0,16,38,1,1,38,4,2,191,1,5,191,2,2,245,1,7,73,1,8,
/* out0295_em-eta15-phi14*/	9,37,0,2,37,1,3,37,2,12,37,3,2,191,2,6,244,2,1,245,0,6,73,0,4,73,1,3,
/* out0296_em-eta16-phi14*/	11,16,4,5,36,2,1,37,0,11,37,3,1,181,2,5,191,2,1,237,1,1,244,2,3,245,0,1,72,2,3,73,0,3,
/* out0297_em-eta17-phi14*/	9,16,4,9,17,0,1,17,1,4,181,1,3,181,2,3,237,1,2,244,2,2,65,1,2,72,2,3,
/* out0298_em-eta18-phi14*/	7,16,1,2,16,2,1,17,0,2,17,1,7,237,1,1,65,1,2,72,2,1,
/* out0299_em-eta19-phi14*/	3,15,3,1,16,0,14,16,1,9,
/* out0300_em-eta0-phi15*/	0,
/* out0301_em-eta1-phi15*/	0,
/* out0302_em-eta2-phi15*/	4,123,1,14,123,2,4,124,1,1,137,2,10,
/* out0303_em-eta3-phi15*/	8,109,1,7,122,0,2,122,1,4,122,2,15,123,0,13,123,1,2,137,0,1,137,2,1,
/* out0304_em-eta4-phi15*/	7,108,0,2,108,1,11,108,2,13,109,0,5,109,1,2,122,0,5,122,2,1,
/* out0305_em-eta5-phi15*/	5,94,1,12,94,2,2,107,2,3,108,0,12,108,2,2,
/* out0306_em-eta6-phi15*/	5,79,1,2,93,2,7,94,0,13,94,1,4,94,2,1,
/* out0307_em-eta7-phi15*/	6,78,1,1,78,2,1,79,0,3,79,1,6,93,0,3,93,2,7,
/* out0308_em-eta8-phi15*/	10,78,0,2,78,1,4,78,2,11,79,0,1,203,1,1,212,1,2,213,0,14,213,1,14,213,2,14,264,1,4,
/* out0309_em-eta9-phi15*/	13,60,1,6,78,0,7,78,2,1,203,0,9,203,1,3,212,1,1,212,2,5,264,0,3,264,1,7,264,2,11,92,0,3,92,1,11,92,2,4,
/* out0310_em-eta10-phi15*/	12,60,0,4,60,1,7,60,2,1,202,1,9,202,2,2,203,0,4,255,1,13,263,2,2,264,2,2,83,1,7,91,2,2,92,2,9,
/* out0311_em-eta11-phi15*/	12,39,4,5,59,2,9,60,0,7,192,1,1,193,0,1,202,2,11,254,2,3,255,0,9,255,1,1,82,2,1,83,0,7,83,1,7,
/* out0312_em-eta12-phi15*/	11,39,4,8,40,1,12,59,2,6,59,3,8,192,0,1,192,1,10,246,1,3,254,2,8,74,1,2,82,2,8,83,0,2,
/* out0313_em-eta13-phi15*/	22,37,5,2,38,2,1,38,5,10,39,0,1,39,1,10,40,1,3,58,3,1,59,3,1,192,0,4,192,2,4,245,1,3,245,2,2,246,0,1,246,1,1,254,0,2,254,2,1,73,1,1,73,2,1,74,0,1,74,1,2,82,0,2,82,2,3,
/* out0314_em-eta14-phi15*/	13,38,2,5,38,3,2,38,4,10,38,5,6,182,0,1,182,1,3,191,2,1,192,0,1,192,2,2,245,1,2,245,2,5,73,1,3,73,2,5,
/* out0315_em-eta15-phi15*/	9,37,2,3,37,3,6,38,3,8,38,4,4,182,0,6,245,0,6,245,2,1,73,0,4,73,2,3,
/* out0316_em-eta16-phi15*/	10,16,4,1,16,5,8,37,3,7,181,2,1,182,0,4,237,1,1,237,2,4,245,0,1,65,2,2,73,0,3,
/* out0317_em-eta17-phi15*/	7,16,5,6,17,0,8,181,1,1,181,2,3,237,1,4,65,1,3,65,2,2,
/* out0318_em-eta18-phi15*/	5,16,2,6,17,0,5,17,4,1,237,1,2,65,1,3,
/* out0319_em-eta19-phi15*/	4,16,0,2,16,1,2,16,2,5,16,3,5,
/* out0320_em-eta0-phi16*/	0,
/* out0321_em-eta1-phi16*/	0,
/* out0322_em-eta2-phi16*/	6,110,1,9,110,2,1,123,2,8,124,0,16,124,1,15,124,2,16,
/* out0323_em-eta3-phi16*/	8,96,1,2,109,1,7,109,2,12,110,0,11,110,1,7,110,2,1,123,0,3,123,2,4,
/* out0324_em-eta4-phi16*/	7,95,1,12,95,2,6,96,0,1,96,1,3,108,2,1,109,0,11,109,2,4,
/* out0325_em-eta5-phi16*/	5,80,1,4,94,2,7,95,0,14,95,1,4,95,2,2,
/* out0326_em-eta6-phi16*/	6,79,1,4,79,2,3,80,0,4,80,1,6,94,0,3,94,2,6,
/* out0327_em-eta7-phi16*/	3,79,0,8,79,1,4,79,2,9,
/* out0328_em-eta8-phi16*/	11,61,1,11,78,2,2,79,0,4,203,1,3,204,0,6,204,1,4,204,2,3,213,0,1,213,1,1,213,2,2,264,1,1,
/* out0329_em-eta9-phi16*/	16,60,2,3,61,0,8,61,1,3,78,2,1,203,0,2,203,1,9,203,2,7,204,0,2,204,1,1,256,0,16,256,1,3,256,2,4,264,1,4,84,0,13,84,1,3,92,1,4,
/* out0330_em-eta10-phi16*/	15,41,1,1,60,0,1,60,2,11,193,0,1,193,1,6,203,0,1,203,2,7,255,1,2,255,2,12,256,2,3,83,1,2,83,2,7,84,0,3,84,2,7,92,1,1,
/* out0331_em-eta11-phi16*/	12,39,4,2,39,5,13,40,5,5,60,0,4,60,2,1,193,0,11,193,1,2,246,1,2,255,0,7,255,2,4,83,0,5,83,2,9,
/* out0332_em-eta12-phi16*/	18,39,2,4,39,4,1,39,5,3,40,0,16,40,1,1,40,4,7,40,5,1,183,0,1,192,1,4,192,2,2,193,0,3,193,2,1,246,0,1,246,1,9,246,2,1,74,1,8,74,2,1,83,0,2,
/* out0333_em-eta13-phi16*/	11,39,0,10,39,1,6,39,2,10,39,3,3,183,0,2,192,2,7,245,2,1,246,0,8,246,1,1,74,0,6,74,1,4,
/* out0334_em-eta14-phi16*/	11,18,4,10,38,2,9,39,0,4,182,1,6,192,2,1,238,1,2,245,2,5,246,0,1,66,1,1,73,2,3,74,0,4,
/* out0335_em-eta15-phi16*/	14,18,1,1,18,4,1,19,1,12,38,2,1,38,3,6,182,0,2,182,1,3,182,2,2,238,0,1,238,1,2,245,0,1,245,2,2,66,1,3,73,2,4,
/* out0336_em-eta16-phi16*/	11,16,5,2,17,5,8,18,1,6,19,1,1,182,0,2,182,2,3,237,2,6,65,2,4,66,0,1,66,1,1,73,0,1,
/* out0337_em-eta17-phi16*/	9,17,4,6,17,5,8,182,0,1,182,2,1,237,0,2,237,1,1,237,2,2,65,0,1,65,2,4,
/* out0338_em-eta18-phi16*/	6,16,2,1,17,3,1,17,4,9,237,1,3,65,0,1,65,1,3,
/* out0339_em-eta19-phi16*/	4,16,2,3,16,3,7,17,3,1,65,1,1,
/* out0340_em-eta0-phi17*/	0,
/* out0341_em-eta1-phi17*/	0,
/* out0342_em-eta2-phi17*/	3,97,0,1,97,1,3,110,2,7,
/* out0343_em-eta3-phi17*/	7,96,1,8,96,2,10,97,0,15,97,1,2,97,2,9,110,0,5,110,2,7,
/* out0344_em-eta4-phi17*/	5,81,1,10,95,2,4,96,0,15,96,1,3,96,2,6,
/* out0345_em-eta5-phi17*/	6,80,1,4,80,2,7,81,0,8,81,1,6,95,0,2,95,2,4,
/* out0346_em-eta6-phi17*/	4,62,1,2,80,0,12,80,1,2,80,2,9,
/* out0347_em-eta7-phi17*/	3,62,0,4,62,1,14,79,2,4,
/* out0348_em-eta8-phi17*/	7,61,1,2,61,2,12,62,0,4,194,1,1,204,0,6,204,1,4,204,2,9,
/* out0349_em-eta9-phi17*/	12,41,1,2,61,0,8,61,2,4,194,0,7,194,1,7,203,2,2,204,0,2,204,1,7,204,2,4,256,1,13,256,2,4,84,1,10,
/* out0350_em-eta10-phi17*/	9,41,0,1,41,1,12,193,1,6,194,0,9,247,1,11,256,2,5,75,1,6,84,1,3,84,2,9,
/* out0351_em-eta11-phi17*/	11,40,2,3,40,5,6,41,0,7,41,1,1,193,1,2,193,2,11,246,2,1,247,0,7,247,1,5,75,0,4,75,1,10,
/* out0352_em-eta12-phi17*/	10,40,2,13,40,3,8,40,4,8,40,5,4,183,1,7,193,2,4,246,2,11,247,0,1,74,2,8,75,0,4,
/* out0353_em-eta13-phi17*/	13,18,5,4,39,0,1,39,2,2,39,3,13,40,3,8,40,4,1,183,0,8,183,1,1,238,1,1,246,0,5,246,2,3,74,0,3,74,2,7,
/* out0354_em-eta14-phi17*/	8,18,4,5,18,5,12,19,0,7,182,1,3,183,0,5,238,1,8,66,1,6,74,0,2,
/* out0355_em-eta15-phi17*/	10,18,1,1,18,2,7,19,0,9,19,1,3,182,1,1,182,2,5,238,0,4,238,1,3,66,0,2,66,1,5,
/* out0356_em-eta16-phi17*/	8,18,0,6,18,1,8,18,2,1,182,2,5,237,2,3,238,0,3,65,2,1,66,0,5,
/* out0357_em-eta17-phi17*/	6,17,2,12,18,0,2,237,0,9,237,2,1,65,0,5,65,2,3,
/* out0358_em-eta18-phi17*/	6,17,2,4,17,3,8,237,0,5,237,1,1,65,0,8,65,1,1,
/* out0359_em-eta19-phi17*/	4,16,3,4,17,3,6,65,0,1,65,1,1,
/* out0360_em-eta0-phi18*/	0,
/* out0361_em-eta1-phi18*/	0,
/* out0362_em-eta2-phi18*/	2,83,1,7,97,1,3,
/* out0363_em-eta3-phi18*/	6,82,1,10,82,2,8,83,0,5,83,1,7,97,1,8,97,2,7,
/* out0364_em-eta4-phi18*/	5,64,1,4,81,2,10,82,0,15,82,1,6,82,2,3,
/* out0365_em-eta5-phi18*/	6,63,1,7,63,2,4,64,0,2,64,1,4,81,0,8,81,2,6,
/* out0366_em-eta6-phi18*/	4,62,2,2,63,0,12,63,1,9,63,2,2,
/* out0367_em-eta7-phi18*/	3,43,1,4,62,0,4,62,2,14,
/* out0368_em-eta8-phi18*/	7,42,1,12,42,2,2,62,0,4,194,1,1,195,0,9,195,1,4,195,2,6,
/* out0369_em-eta9-phi18*/	14,41,2,2,42,0,8,42,1,4,185,0,2,194,1,7,194,2,7,195,0,4,195,1,7,195,2,2,248,0,16,248,1,6,248,2,5,76,0,10,76,1,6,
/* out0370_em-eta10-phi18*/	9,41,0,1,41,2,12,184,1,6,194,2,9,247,2,11,248,2,5,75,2,6,76,0,6,76,2,10,
/* out0371_em-eta11-phi18*/	11,20,4,3,20,5,6,41,0,7,41,2,1,184,0,11,184,1,2,239,1,1,247,0,7,247,2,5,75,0,4,75,2,10,
/* out0372_em-eta12-phi18*/	10,20,4,13,20,5,4,21,0,8,21,1,8,183,1,7,184,0,4,239,1,11,247,0,1,67,1,8,75,0,4,
/* out0373_em-eta13-phi18*/	13,19,5,4,20,0,1,20,1,13,20,2,2,21,0,1,21,1,8,183,1,1,183,2,8,238,2,1,239,0,5,239,1,3,67,0,3,67,1,7,
/* out0374_em-eta14-phi18*/	8,19,2,5,19,4,7,19,5,12,177,1,3,183,2,5,238,2,8,66,2,6,67,0,2,
/* out0375_em-eta15-phi18*/	10,18,2,7,18,3,1,19,3,3,19,4,9,177,0,5,177,1,1,238,0,4,238,2,3,66,0,2,66,2,5,
/* out0376_em-eta16-phi18*/	8,18,0,6,18,2,1,18,3,8,177,0,5,232,2,3,238,0,3,60,2,1,66,0,5,
/* out0377_em-eta17-phi18*/	5,0,4,12,18,0,2,232,1,4,60,1,2,60,2,2,
/* out0378_em-eta18-phi18*/	4,0,4,4,1,1,8,232,1,3,60,1,3,
/* out0379_em-eta19-phi18*/	3,0,1,4,1,1,6,60,1,1,
/* out0380_em-eta0-phi19*/	0,
/* out0381_em-eta1-phi19*/	0,
/* out0382_em-eta2-phi19*/	6,66,1,8,83,1,1,83,2,9,84,0,16,84,1,16,84,2,15,
/* out0383_em-eta3-phi19*/	8,65,1,12,65,2,7,66,0,3,66,1,4,82,2,2,83,0,11,83,1,1,83,2,7,
/* out0384_em-eta4-phi19*/	7,45,1,1,64,1,6,64,2,12,65,0,11,65,1,4,82,0,1,82,2,3,
/* out0385_em-eta5-phi19*/	5,44,1,7,63,2,4,64,0,14,64,1,2,64,2,4,
/* out0386_em-eta6-phi19*/	6,43,1,3,43,2,4,44,0,3,44,1,6,63,0,4,63,2,6,
/* out0387_em-eta7-phi19*/	3,43,0,8,43,1,9,43,2,4,
/* out0388_em-eta8-phi19*/	12,23,1,2,42,2,11,43,0,4,185,1,3,186,0,2,186,1,1,186,2,1,195,0,3,195,1,4,195,2,6,241,1,1,248,1,1,
/* out0389_em-eta9-phi19*/	16,22,1,3,23,1,1,42,0,8,42,2,3,185,0,7,185,1,9,185,2,2,195,1,1,195,2,2,241,0,10,241,2,1,248,1,9,248,2,3,69,0,8,69,1,1,76,1,8,
/* out0390_em-eta10-phi19*/	16,22,0,1,22,1,11,41,2,1,184,1,6,184,2,1,185,0,7,185,2,1,240,1,12,240,2,2,248,2,3,68,1,7,68,2,2,69,0,2,69,2,1,76,1,2,76,2,6,
/* out0391_em-eta11-phi19*/	12,20,5,5,21,2,2,21,5,13,22,0,4,22,1,1,184,1,2,184,2,11,239,2,2,240,0,7,240,1,4,68,0,5,68,1,9,
/* out0392_em-eta12-phi19*/	18,20,2,4,20,5,1,21,0,7,21,2,1,21,3,1,21,4,16,21,5,3,178,0,2,178,1,4,183,2,1,184,0,1,184,2,3,239,0,1,239,1,1,239,2,9,67,1,1,67,2,8,68,0,2,
/* out0393_em-eta13-phi19*/	11,20,0,10,20,1,3,20,2,10,20,3,6,178,0,7,183,2,2,233,1,1,239,0,8,239,2,1,67,0,6,67,2,4,
/* out0394_em-eta14-phi19*/	11,2,4,9,19,2,10,20,0,4,177,1,6,178,0,1,233,1,5,238,2,2,239,0,1,61,1,3,66,2,1,67,0,4,
/* out0395_em-eta15-phi19*/	14,2,4,1,3,1,6,18,3,1,19,2,1,19,3,12,177,0,2,177,1,3,177,2,2,233,0,1,233,1,2,238,0,1,238,2,2,61,1,4,66,2,3,
/* out0396_em-eta16-phi19*/	11,0,5,8,1,5,2,18,3,6,19,3,1,177,0,3,177,2,2,232,2,6,60,2,4,61,0,1,66,0,1,66,2,1,
/* out0397_em-eta17-phi19*/	8,0,5,8,1,0,6,177,0,1,177,2,1,232,1,2,232,2,2,60,1,1,60,2,4,
/* out0398_em-eta18-phi19*/	5,0,2,1,1,0,9,1,1,1,232,1,3,60,1,4,
/* out0399_em-eta19-phi19*/	4,0,1,7,0,2,3,1,1,1,60,1,1,
/* out0400_em-eta0-phi20*/	0,
/* out0401_em-eta1-phi20*/	0,
/* out0402_em-eta2-phi20*/	4,47,1,10,66,1,4,66,2,14,84,2,1,
/* out0403_em-eta3-phi20*/	8,46,0,2,46,1,15,46,2,4,47,0,1,47,1,1,65,2,7,66,0,13,66,2,2,
/* out0404_em-eta4-phi20*/	7,45,0,2,45,1,13,45,2,11,46,0,5,46,1,1,65,0,5,65,2,2,
/* out0405_em-eta5-phi20*/	5,25,1,3,44,1,2,44,2,12,45,0,12,45,1,2,
/* out0406_em-eta6-phi20*/	5,24,1,7,43,2,2,44,0,13,44,1,1,44,2,4,
/* out0407_em-eta7-phi20*/	6,23,1,1,23,2,1,24,0,3,24,1,7,43,0,3,43,2,6,
/* out0408_em-eta8-phi20*/	10,23,0,2,23,1,11,23,2,4,43,0,1,180,1,2,185,1,1,186,0,14,186,1,14,186,2,14,241,1,4,
/* out0409_em-eta9-phi20*/	13,22,2,6,23,0,7,23,1,1,180,0,5,180,1,1,185,1,3,185,2,9,241,0,6,241,1,6,241,2,11,69,0,6,69,1,10,69,2,4,
/* out0410_em-eta10-phi20*/	12,22,0,4,22,1,1,22,2,7,179,0,2,179,1,9,185,2,4,235,1,2,240,2,13,241,2,1,63,1,2,68,2,7,69,2,9,
/* out0411_em-eta11-phi20*/	12,4,4,9,21,2,5,22,0,7,178,1,1,179,0,11,184,2,1,234,1,3,240,0,9,240,2,1,62,1,1,68,0,7,68,2,7,
/* out0412_em-eta12-phi20*/	11,4,4,6,5,1,8,21,2,8,21,3,12,178,1,10,178,2,1,234,1,8,239,2,3,62,1,8,67,2,2,68,0,2,
/* out0413_em-eta13-phi20*/	22,2,4,1,2,5,10,3,5,2,4,1,1,5,1,1,20,0,1,20,3,10,21,3,3,178,0,4,178,2,4,233,1,2,233,2,3,234,0,2,234,1,1,239,0,1,239,2,1,61,1,1,61,2,1,62,0,2,62,1,3,67,0,1,67,2,2,
/* out0414_em-eta14-phi20*/	13,2,4,5,2,5,6,3,0,10,3,1,2,173,0,1,177,1,3,177,2,1,178,0,2,178,2,1,233,1,5,233,2,2,61,1,5,61,2,3,
/* out0415_em-eta15-phi20*/	9,2,1,6,2,2,3,3,0,4,3,1,8,177,2,6,233,0,6,233,1,1,61,0,4,61,1,3,
/* out0416_em-eta16-phi20*/	10,1,2,1,1,5,8,2,1,7,172,1,1,177,2,4,232,0,1,232,2,4,233,0,1,60,2,2,61,0,3,
/* out0417_em-eta17-phi20*/	8,1,4,8,1,5,6,172,1,4,232,0,6,232,1,1,232,2,1,60,0,6,60,2,3,
/* out0418_em-eta18-phi20*/	6,0,2,6,1,0,1,1,4,5,232,1,2,60,0,1,60,1,3,
/* out0419_em-eta19-phi20*/	4,0,0,2,0,1,5,0,2,5,0,3,2,
/* out0420_em-eta0-phi21*/	0,
/* out0421_em-eta1-phi21*/	0,
/* out0422_em-eta2-phi21*/	7,27,1,1,27,2,1,28,0,9,28,2,1,47,0,7,47,1,5,47,2,16,
/* out0423_em-eta3-phi21*/	7,26,2,1,27,0,4,27,1,15,27,2,1,46,0,4,46,2,12,47,0,8,
/* out0424_em-eta4-phi21*/	5,26,0,7,26,1,16,26,2,6,45,2,5,46,0,5,
/* out0425_em-eta5-phi21*/	5,25,0,4,25,1,12,25,2,12,26,0,2,45,0,2,
/* out0426_em-eta6-phi21*/	5,8,1,2,24,1,1,24,2,12,25,0,10,25,1,1,
/* out0427_em-eta7-phi21*/	5,7,1,3,23,2,1,24,0,13,24,1,1,24,2,4,
/* out0428_em-eta8-phi21*/	9,7,1,5,23,0,2,23,2,10,180,1,10,180,2,1,186,1,1,186,2,1,236,0,7,241,1,2,
/* out0429_em-eta9-phi21*/	17,6,1,9,6,2,1,23,0,5,180,0,9,180,1,3,180,2,7,235,1,3,235,2,3,236,0,5,236,2,3,241,1,3,241,2,3,63,2,1,64,0,12,64,2,3,69,1,5,69,2,1,
/* out0430_em-eta10-phi21*/	16,4,5,1,5,5,1,6,0,3,6,1,6,22,2,3,175,0,1,179,1,7,179,2,6,180,0,2,235,0,4,235,1,10,235,2,2,63,0,1,63,1,11,63,2,5,69,2,1,
/* out0431_em-eta11-phi21*/	16,4,4,1,4,5,15,5,0,6,5,4,6,5,5,11,174,1,1,179,0,2,179,2,9,234,1,2,234,2,7,235,0,4,235,1,1,62,1,1,62,2,3,63,0,7,63,1,3,
/* out0432_em-eta12-phi21*/	16,4,1,6,4,2,9,5,0,10,5,1,7,5,4,1,174,0,4,174,1,2,178,1,1,178,2,4,179,0,1,234,0,5,234,1,2,234,2,3,62,0,1,62,1,3,62,2,7,
/* out0433_em-eta13-phi21*/	11,3,2,5,3,5,11,4,0,4,4,1,9,173,1,2,174,0,1,178,2,6,229,1,1,233,2,3,234,0,6,62,0,10,
/* out0434_em-eta14-phi21*/	10,2,2,1,3,0,2,3,2,1,3,3,1,3,4,16,3,5,3,173,0,2,173,1,5,233,2,7,61,2,8,
/* out0435_em-eta15-phi21*/	9,2,0,2,2,1,2,2,2,12,2,3,3,173,0,6,228,1,1,233,0,6,61,0,4,61,2,3,
/* out0436_em-eta16-phi21*/	11,1,2,5,2,0,11,2,1,1,172,1,2,172,2,3,173,0,1,228,1,3,232,0,2,233,0,1,56,1,3,61,0,3,
/* out0437_em-eta17-phi21*/	9,1,2,9,1,3,4,1,4,1,172,1,5,172,2,1,228,1,2,232,0,6,56,1,3,60,0,5,
/* out0438_em-eta18-phi21*/	11,0,2,1,0,3,2,1,3,7,1,4,2,228,0,1,232,0,1,232,1,1,56,0,2,56,1,1,60,0,4,60,1,1,
/* out0439_em-eta19-phi21*/	2,0,0,14,0,3,9,
/* out0440_em-eta0-phi22*/	0,
/* out0441_em-eta1-phi22*/	0,
/* out0442_em-eta2-phi22*/	5,11,1,8,11,2,2,27,2,1,28,0,7,28,2,15,
/* out0443_em-eta3-phi22*/	6,10,1,7,10,2,4,11,0,3,11,1,8,27,0,12,27,2,13,
/* out0444_em-eta4-phi22*/	6,9,1,3,9,2,5,10,0,6,10,1,9,26,0,6,26,2,9,
/* out0445_em-eta5-phi22*/	7,8,2,2,9,0,8,9,1,13,9,2,2,25,0,1,25,2,4,26,0,1,
/* out0446_em-eta6-phi22*/	4,8,0,4,8,1,13,8,2,8,25,0,1,
/* out0447_em-eta7-phi22*/	4,7,1,4,7,2,10,8,0,6,8,1,1,
/* out0448_em-eta8-phi22*/	7,7,0,12,7,1,4,7,2,2,176,0,8,180,2,2,236,0,4,236,2,1,
/* out0449_em-eta9-phi22*/	13,6,1,1,6,2,13,7,0,1,175,1,7,176,0,4,176,2,3,180,2,6,231,1,7,235,2,4,236,2,12,59,1,3,64,0,4,64,2,13,
/* out0450_em-eta10-phi22*/	14,6,0,11,175,0,9,175,1,6,230,1,1,230,2,3,231,0,1,231,1,2,235,0,5,235,2,7,58,2,1,59,0,3,59,1,5,63,0,1,63,2,10,
/* out0451_em-eta11-phi22*/	14,5,2,16,5,3,8,5,4,5,5,5,4,174,1,8,175,0,4,179,2,1,230,1,9,234,2,2,235,0,3,58,1,7,58,2,1,62,2,1,63,0,7,
/* out0452_em-eta12-phi22*/	17,4,0,2,4,2,7,4,3,14,5,3,6,5,4,4,174,0,5,174,1,3,174,2,2,229,1,1,229,2,1,230,0,1,230,1,3,234,0,2,234,2,4,58,0,1,58,1,6,62,2,5,
/* out0453_em-eta13-phi22*/	11,3,2,5,4,0,10,173,1,4,174,0,5,229,1,8,229,2,3,234,0,1,57,1,6,57,2,2,58,0,1,62,0,3,
/* out0454_em-eta14-phi22*/	9,3,2,5,3,3,13,173,1,5,173,2,2,229,0,2,229,1,5,233,2,1,57,0,1,57,1,8,
/* out0455_em-eta15-phi22*/	15,2,0,1,2,3,13,3,3,2,173,0,4,173,2,3,228,1,3,228,2,3,229,0,1,233,0,1,56,1,1,56,2,2,57,0,2,57,1,1,61,0,1,61,2,1,
/* out0456_em-eta16-phi22*/	8,2,0,2,172,2,4,173,0,2,228,0,1,228,1,5,228,2,1,56,1,4,56,2,4,
/* out0457_em-eta17-phi22*/	7,1,2,1,172,1,2,172,2,4,228,0,3,228,1,2,56,0,2,56,1,4,
/* out0458_em-eta18-phi22*/	4,1,3,5,172,1,1,228,0,2,56,0,3,
/* out0459_em-eta19-phi22*/	1,0,3,3,
/* out0460_em-eta0-phi23*/	0,
/* out0461_em-eta1-phi23*/	0,
/* out0462_em-eta2-phi23*/	1,11,2,13,
/* out0463_em-eta3-phi23*/	3,10,2,9,11,0,13,11,2,1,
/* out0464_em-eta4-phi23*/	3,9,2,4,10,0,10,10,2,3,
/* out0465_em-eta5-phi23*/	2,9,0,8,9,2,5,
/* out0466_em-eta6-phi23*/	2,8,0,4,8,2,6,
/* out0467_em-eta7-phi23*/	2,7,2,2,8,0,2,
/* out0468_em-eta8-phi23*/	5,7,0,3,7,2,2,176,0,4,176,2,4,231,2,2,
/* out0469_em-eta9-phi23*/	9,6,2,2,175,1,3,175,2,3,176,2,9,231,0,3,231,1,6,231,2,14,59,1,4,59,2,11,
/* out0470_em-eta10-phi23*/	10,6,0,2,175,0,1,175,2,12,230,2,6,231,0,12,231,1,1,58,2,1,59,0,12,59,1,4,59,2,5,
/* out0471_em-eta11-phi23*/	11,174,1,2,174,2,3,175,0,1,175,2,1,230,0,4,230,1,3,230,2,7,58,0,2,58,1,2,58,2,12,59,0,1,
/* out0472_em-eta12-phi23*/	8,4,3,2,5,3,2,174,2,9,229,2,4,230,0,11,58,0,11,58,1,1,58,2,1,
/* out0473_em-eta13-phi23*/	8,173,2,1,174,0,1,174,2,2,229,0,1,229,1,1,229,2,8,57,2,12,58,0,1,
/* out0474_em-eta14-phi23*/	5,173,2,5,229,0,8,57,0,6,57,1,1,57,2,2,
/* out0475_em-eta15-phi23*/	5,173,2,4,228,2,8,229,0,4,56,2,3,57,0,7,
/* out0476_em-eta16-phi23*/	5,172,2,1,173,2,1,228,0,2,228,2,4,56,2,6,
/* out0477_em-eta17-phi23*/	4,172,2,3,228,0,5,56,0,5,56,2,1,
/* out0478_em-eta18-phi23*/	3,172,1,1,228,0,2,56,0,4,
/* out0479_em-eta19-phi23*/	0
};