parameter integer matrixH [0:5880] = {
/* num inputs = 158(in0-in157) */
/* num outputs = 480(out0-out479) */
//* max inputs per outputs = 9 */
//* total number of input in adders 1800 */

/* out0000_had-eta0-phi0*/	1, 113, 0, 4, 
/* out0001_had-eta1-phi0*/	1, 113, 0, 4, 
/* out0002_had-eta2-phi0*/	1, 112, 0, 4, 
/* out0003_had-eta3-phi0*/	4, 35, 2, 6, 36, 1, 10, 111, 0, 1, 112, 0, 4, 
/* out0004_had-eta4-phi0*/	7, 27, 0, 11, 27, 1, 12, 27, 2, 16, 34, 2, 1, 35, 1, 8, 35, 2, 3, 111, 0, 4, 
/* out0005_had-eta5-phi0*/	8, 26, 0, 3, 26, 2, 15, 27, 0, 5, 27, 1, 4, 34, 1, 4, 34, 2, 5, 110, 0, 1, 111, 0, 3, 
/* out0006_had-eta6-phi0*/	6, 26, 0, 13, 26, 1, 15, 26, 2, 1, 33, 2, 4, 34, 1, 1, 110, 0, 3, 
/* out0007_had-eta7-phi0*/	7, 25, 0, 9, 25, 1, 11, 25, 2, 16, 26, 1, 1, 33, 1, 3, 33, 2, 1, 110, 0, 3, 
/* out0008_had-eta8-phi0*/	5, 24, 2, 12, 25, 0, 7, 25, 1, 5, 32, 2, 2, 110, 0, 1, 
/* out0009_had-eta9-phi0*/	4, 24, 0, 8, 24, 1, 11, 24, 2, 4, 32, 1, 1, 
/* out0010_had-eta10-phi0*/	3, 5, 11, 1, 24, 0, 6, 24, 1, 4, 
/* out0011_had-eta11-phi0*/	8, 3, 2, 1, 3, 3, 11, 3, 8, 16, 3, 9, 16, 3, 10, 3, 5, 5, 2, 5, 11, 1, 24, 1, 1, 
/* out0012_had-eta12-phi0*/	6, 3, 0, 1, 3, 1, 4, 3, 2, 15, 3, 3, 3, 3, 6, 14, 3, 10, 13, 
/* out0013_had-eta13-phi0*/	6, 1, 8, 1, 1, 9, 4, 3, 1, 7, 3, 4, 16, 3, 6, 2, 3, 7, 16, 
/* out0014_had-eta14-phi0*/	5, 1, 2, 1, 1, 3, 6, 1, 8, 15, 1, 9, 12, 1, 10, 2, 
/* out0015_had-eta15-phi0*/	4, 1, 2, 12, 1, 3, 1, 1, 6, 12, 1, 10, 14, 
/* out0016_had-eta16-phi0*/	4, 1, 1, 3, 1, 2, 3, 1, 6, 4, 1, 7, 4, 
/* out0017_had-eta17-phi0*/	4, 0, 3, 16, 0, 4, 4, 1, 4, 16, 1, 7, 11, 
/* out0018_had-eta18-phi0*/	4, 0, 1, 1, 0, 2, 1, 0, 4, 10, 0, 5, 11, 
/* out0019_had-eta19-phi0*/	2, 0, 1, 13, 0, 5, 5, 
/* out0020_had-eta0-phi1*/	1, 113, 0, 4, 
/* out0021_had-eta1-phi1*/	1, 113, 0, 4, 
/* out0022_had-eta2-phi1*/	3, 36, 0, 3, 46, 2, 1, 112, 0, 4, 
/* out0023_had-eta3-phi1*/	8, 35, 0, 6, 35, 2, 6, 36, 0, 13, 36, 1, 6, 46, 1, 7, 46, 2, 8, 111, 0, 1, 112, 0, 4, 
/* out0024_had-eta4-phi1*/	8, 34, 0, 1, 34, 2, 4, 35, 0, 10, 35, 1, 8, 35, 2, 1, 45, 1, 2, 45, 2, 4, 111, 0, 4, 
/* out0025_had-eta5-phi1*/	5, 34, 0, 13, 34, 1, 7, 34, 2, 6, 110, 0, 1, 111, 0, 3, 
/* out0026_had-eta6-phi1*/	4, 33, 0, 5, 33, 2, 11, 34, 1, 4, 110, 0, 3, 
/* out0027_had-eta7-phi1*/	4, 32, 2, 2, 33, 0, 3, 33, 1, 13, 110, 0, 3, 
/* out0028_had-eta8-phi1*/	4, 32, 0, 1, 32, 1, 2, 32, 2, 11, 110, 0, 1, 
/* out0029_had-eta9-phi1*/	4, 5, 8, 4, 5, 9, 1, 24, 0, 1, 32, 1, 10, 
/* out0030_had-eta10-phi1*/	5, 5, 8, 12, 5, 9, 3, 5, 10, 9, 5, 11, 12, 24, 0, 1, 
/* out0031_had-eta11-phi1*/	6, 3, 0, 2, 3, 3, 2, 5, 4, 7, 5, 5, 14, 5, 6, 7, 5, 11, 2, 
/* out0032_had-eta12-phi1*/	4, 3, 0, 13, 3, 1, 1, 4, 8, 9, 5, 4, 5, 
/* out0033_had-eta13-phi1*/	5, 3, 1, 4, 4, 5, 3, 4, 8, 1, 4, 10, 1, 4, 11, 15, 
/* out0034_had-eta14-phi1*/	4, 1, 0, 1, 1, 3, 6, 4, 4, 2, 4, 5, 10, 
/* out0035_had-eta15-phi1*/	4, 1, 0, 12, 1, 1, 1, 1, 3, 3, 4, 4, 1, 
/* out0036_had-eta16-phi1*/	4, 1, 0, 2, 1, 1, 9, 2, 8, 1, 2, 11, 2, 
/* out0037_had-eta17-phi1*/	6, 0, 2, 1, 0, 4, 1, 1, 1, 3, 1, 7, 1, 2, 5, 2, 2, 11, 4, 
/* out0038_had-eta18-phi1*/	3, 0, 2, 9, 0, 4, 1, 2, 5, 1, 
/* out0039_had-eta19-phi1*/	3, 0, 0, 1, 0, 1, 2, 0, 2, 4, 
/* out0040_had-eta0-phi2*/	1, 117, 0, 4, 
/* out0041_had-eta1-phi2*/	1, 117, 0, 4, 
/* out0042_had-eta2-phi2*/	3, 46, 0, 1, 46, 2, 3, 116, 0, 4, 
/* out0043_had-eta3-phi2*/	8, 45, 2, 1, 46, 0, 15, 46, 1, 9, 46, 2, 4, 55, 1, 1, 55, 2, 5, 115, 0, 1, 116, 0, 4, 
/* out0044_had-eta4-phi2*/	5, 45, 0, 12, 45, 1, 7, 45, 2, 11, 55, 1, 1, 115, 0, 4, 
/* out0045_had-eta5-phi2*/	7, 34, 0, 2, 44, 0, 2, 44, 2, 15, 45, 0, 1, 45, 1, 7, 114, 0, 1, 115, 0, 3, 
/* out0046_had-eta6-phi2*/	5, 33, 0, 4, 43, 2, 2, 44, 1, 13, 44, 2, 1, 114, 0, 3, 
/* out0047_had-eta7-phi2*/	5, 32, 2, 1, 33, 0, 4, 43, 1, 4, 43, 2, 8, 114, 0, 3, 
/* out0048_had-eta8-phi2*/	4, 32, 0, 11, 42, 2, 1, 43, 1, 3, 114, 0, 1, 
/* out0049_had-eta9-phi2*/	6, 5, 3, 3, 5, 9, 6, 32, 0, 4, 32, 1, 3, 42, 1, 1, 42, 2, 2, 
/* out0050_had-eta10-phi2*/	6, 5, 0, 1, 5, 1, 1, 5, 2, 11, 5, 3, 13, 5, 9, 6, 5, 10, 7, 
/* out0051_had-eta11-phi2*/	5, 5, 1, 6, 5, 2, 5, 5, 4, 1, 5, 6, 9, 5, 7, 12, 
/* out0052_had-eta12-phi2*/	5, 4, 8, 6, 4, 9, 14, 4, 10, 2, 5, 4, 3, 5, 7, 3, 
/* out0053_had-eta13-phi2*/	4, 4, 2, 2, 4, 6, 7, 4, 10, 13, 4, 11, 1, 
/* out0054_had-eta14-phi2*/	4, 4, 4, 6, 4, 5, 3, 4, 6, 7, 4, 7, 3, 
/* out0055_had-eta15-phi2*/	3, 1, 0, 1, 2, 8, 9, 4, 4, 7, 
/* out0056_had-eta16-phi2*/	3, 2, 8, 5, 2, 10, 2, 2, 11, 6, 
/* out0057_had-eta17-phi2*/	4, 2, 5, 5, 2, 6, 1, 2, 10, 1, 2, 11, 4, 
/* out0058_had-eta18-phi2*/	4, 0, 0, 3, 0, 2, 1, 2, 4, 3, 2, 5, 6, 
/* out0059_had-eta19-phi2*/	2, 0, 0, 12, 2, 4, 1, 
/* out0060_had-eta0-phi3*/	1, 117, 0, 4, 
/* out0061_had-eta1-phi3*/	1, 117, 0, 4, 
/* out0062_had-eta2-phi3*/	1, 116, 0, 4, 
/* out0063_had-eta3-phi3*/	6, 55, 0, 14, 55, 1, 5, 55, 2, 11, 104, 1, 5, 115, 0, 1, 116, 0, 4, 
/* out0064_had-eta4-phi3*/	6, 45, 0, 3, 54, 0, 3, 54, 2, 15, 55, 0, 1, 55, 1, 9, 115, 0, 4, 
/* out0065_had-eta5-phi3*/	6, 44, 0, 9, 53, 2, 3, 54, 1, 13, 54, 2, 1, 114, 0, 1, 115, 0, 3, 
/* out0066_had-eta6-phi3*/	7, 43, 0, 2, 43, 2, 3, 44, 0, 5, 44, 1, 3, 53, 1, 3, 53, 2, 5, 114, 0, 3, 
/* out0067_had-eta7-phi3*/	4, 43, 0, 11, 43, 1, 3, 43, 2, 3, 114, 0, 3, 
/* out0068_had-eta8-phi3*/	4, 42, 2, 8, 43, 0, 1, 43, 1, 6, 114, 0, 1, 
/* out0069_had-eta9-phi3*/	3, 42, 0, 1, 42, 1, 6, 42, 2, 5, 
/* out0070_had-eta10-phi3*/	3, 5, 0, 13, 6, 8, 9, 42, 1, 5, 
/* out0071_had-eta11-phi3*/	6, 5, 0, 2, 5, 1, 9, 5, 7, 1, 6, 5, 3, 6, 8, 4, 6, 11, 15, 
/* out0072_had-eta12-phi3*/	6, 4, 0, 3, 4, 2, 1, 4, 3, 14, 4, 9, 2, 6, 4, 1, 6, 5, 8, 
/* out0073_had-eta13-phi3*/	4, 4, 0, 4, 4, 1, 5, 4, 2, 12, 4, 3, 2, 
/* out0074_had-eta14-phi3*/	4, 4, 1, 6, 4, 2, 1, 4, 6, 2, 4, 7, 11, 
/* out0075_had-eta15-phi3*/	3, 2, 8, 1, 2, 9, 13, 4, 7, 2, 
/* out0076_had-eta16-phi3*/	3, 2, 2, 1, 2, 9, 2, 2, 10, 11, 
/* out0077_had-eta17-phi3*/	2, 2, 6, 9, 2, 10, 2, 
/* out0078_had-eta18-phi3*/	4, 2, 4, 5, 2, 5, 2, 2, 6, 2, 2, 7, 1, 
/* out0079_had-eta19-phi3*/	1, 2, 4, 5, 
/* out0080_had-eta0-phi4*/	1, 121, 0, 4, 
/* out0081_had-eta1-phi4*/	1, 121, 0, 4, 
/* out0082_had-eta2-phi4*/	4, 104, 0, 12, 104, 1, 1, 105, 1, 5, 120, 0, 4, 
/* out0083_had-eta3-phi4*/	9, 55, 0, 1, 103, 0, 7, 103, 2, 14, 104, 0, 4, 104, 1, 10, 105, 0, 1, 105, 1, 4, 119, 0, 1, 120, 0, 4, 
/* out0084_had-eta4-phi4*/	5, 54, 0, 9, 102, 2, 6, 103, 1, 14, 103, 2, 2, 119, 0, 4, 
/* out0085_had-eta5-phi4*/	8, 53, 0, 5, 53, 2, 5, 54, 0, 4, 54, 1, 3, 102, 1, 4, 102, 2, 4, 118, 0, 1, 119, 0, 3, 
/* out0086_had-eta6-phi4*/	4, 53, 0, 7, 53, 1, 11, 53, 2, 3, 118, 0, 3, 
/* out0087_had-eta7-phi4*/	4, 43, 0, 2, 52, 2, 14, 53, 1, 2, 118, 0, 3, 
/* out0088_had-eta8-phi4*/	4, 42, 0, 6, 52, 1, 8, 52, 2, 1, 118, 0, 1, 
/* out0089_had-eta9-phi4*/	3, 42, 0, 9, 42, 1, 2, 60, 2, 1, 
/* out0090_had-eta10-phi4*/	6, 6, 2, 1, 6, 3, 6, 6, 8, 3, 6, 9, 16, 6, 10, 2, 42, 1, 2, 
/* out0091_had-eta11-phi4*/	4, 6, 2, 7, 6, 6, 11, 6, 10, 14, 6, 11, 1, 
/* out0092_had-eta12-phi4*/	5, 4, 0, 1, 6, 4, 14, 6, 5, 5, 6, 6, 4, 6, 7, 3, 
/* out0093_had-eta13-phi4*/	4, 4, 0, 8, 4, 1, 1, 7, 8, 10, 7, 11, 2, 
/* out0094_had-eta14-phi4*/	3, 4, 1, 4, 7, 5, 3, 7, 11, 10, 
/* out0095_had-eta15-phi4*/	3, 2, 3, 12, 2, 9, 1, 7, 5, 2, 
/* out0096_had-eta16-phi4*/	2, 2, 2, 9, 2, 3, 4, 
/* out0097_had-eta17-phi4*/	3, 2, 1, 2, 2, 2, 6, 2, 6, 4, 
/* out0098_had-eta18-phi4*/	1, 2, 7, 9, 
/* out0099_had-eta19-phi4*/	2, 2, 4, 2, 2, 7, 1, 
/* out0100_had-eta0-phi5*/	1, 121, 0, 4, 
/* out0101_had-eta1-phi5*/	1, 121, 0, 4, 
/* out0102_had-eta2-phi5*/	2, 105, 1, 4, 120, 0, 4, 
/* out0103_had-eta3-phi5*/	6, 92, 2, 12, 103, 0, 6, 105, 0, 15, 105, 1, 3, 119, 0, 1, 120, 0, 4, 
/* out0104_had-eta4-phi5*/	7, 92, 1, 8, 92, 2, 4, 102, 0, 10, 102, 2, 5, 103, 0, 3, 103, 1, 2, 119, 0, 4, 
/* out0105_had-eta5-phi5*/	7, 53, 0, 1, 90, 2, 5, 102, 0, 6, 102, 1, 12, 102, 2, 1, 118, 0, 1, 119, 0, 3, 
/* out0106_had-eta6-phi5*/	4, 53, 0, 3, 90, 1, 6, 90, 2, 11, 118, 0, 3, 
/* out0107_had-eta7-phi5*/	5, 52, 0, 14, 52, 1, 1, 52, 2, 1, 90, 1, 2, 118, 0, 3, 
/* out0108_had-eta8-phi5*/	4, 52, 0, 2, 52, 1, 7, 60, 2, 5, 118, 0, 1, 
/* out0109_had-eta9-phi5*/	2, 60, 1, 2, 60, 2, 10, 
/* out0110_had-eta10-phi5*/	3, 6, 0, 7, 6, 3, 9, 60, 1, 6, 
/* out0111_had-eta11-phi5*/	5, 6, 0, 9, 6, 1, 13, 6, 2, 8, 6, 3, 1, 6, 6, 1, 
/* out0112_had-eta12-phi5*/	5, 6, 1, 3, 6, 4, 1, 6, 7, 13, 7, 8, 2, 7, 9, 8, 
/* out0113_had-eta13-phi5*/	4, 7, 8, 4, 7, 9, 7, 7, 10, 10, 7, 11, 2, 
/* out0114_had-eta14-phi5*/	4, 7, 5, 5, 7, 6, 7, 7, 10, 5, 7, 11, 2, 
/* out0115_had-eta15-phi5*/	3, 2, 0, 3, 7, 4, 7, 7, 5, 6, 
/* out0116_had-eta16-phi5*/	2, 2, 0, 12, 2, 1, 1, 
/* out0117_had-eta17-phi5*/	2, 2, 0, 1, 2, 1, 10, 
/* out0118_had-eta18-phi5*/	2, 2, 1, 3, 2, 7, 5, 
/* out0119_had-eta19-phi5*/	0, 
/* out0120_had-eta0-phi6*/	1, 125, 0, 4, 
/* out0121_had-eta1-phi6*/	1, 125, 0, 4, 
/* out0122_had-eta2-phi6*/	2, 94, 0, 4, 124, 0, 4, 
/* out0123_had-eta3-phi6*/	6, 92, 0, 12, 93, 2, 6, 94, 0, 3, 94, 1, 15, 123, 0, 1, 124, 0, 4, 
/* out0124_had-eta4-phi6*/	7, 91, 0, 5, 91, 2, 10, 92, 0, 4, 92, 1, 8, 93, 1, 2, 93, 2, 3, 123, 0, 4, 
/* out0125_had-eta5-phi6*/	7, 62, 2, 1, 90, 0, 5, 91, 0, 1, 91, 1, 12, 91, 2, 6, 122, 0, 1, 123, 0, 3, 
/* out0126_had-eta6-phi6*/	4, 62, 2, 3, 90, 0, 11, 90, 1, 6, 122, 0, 3, 
/* out0127_had-eta7-phi6*/	5, 61, 0, 1, 61, 1, 1, 61, 2, 14, 90, 1, 2, 122, 0, 3, 
/* out0128_had-eta8-phi6*/	4, 60, 0, 5, 61, 1, 7, 61, 2, 2, 122, 0, 1, 
/* out0129_had-eta9-phi6*/	2, 60, 0, 10, 60, 1, 2, 
/* out0130_had-eta10-phi6*/	3, 8, 8, 7, 8, 9, 9, 60, 1, 6, 
/* out0131_had-eta11-phi6*/	5, 8, 6, 1, 8, 8, 9, 8, 9, 1, 8, 10, 8, 8, 11, 13, 
/* out0132_had-eta12-phi6*/	6, 7, 0, 1, 7, 3, 9, 7, 9, 1, 8, 4, 1, 8, 5, 13, 8, 11, 3, 
/* out0133_had-eta13-phi6*/	5, 7, 0, 3, 7, 1, 1, 7, 2, 11, 7, 3, 7, 7, 10, 1, 
/* out0134_had-eta14-phi6*/	4, 7, 1, 1, 7, 2, 5, 7, 6, 9, 7, 7, 4, 
/* out0135_had-eta15-phi6*/	3, 7, 4, 9, 7, 7, 5, 9, 8, 3, 
/* out0136_had-eta16-phi6*/	2, 9, 8, 12, 9, 11, 1, 
/* out0137_had-eta17-phi6*/	2, 9, 8, 1, 9, 11, 10, 
/* out0138_had-eta18-phi6*/	2, 9, 5, 5, 9, 11, 3, 
/* out0139_had-eta19-phi6*/	0, 
/* out0140_had-eta0-phi7*/	1, 125, 0, 4, 
/* out0141_had-eta1-phi7*/	1, 125, 0, 4, 
/* out0142_had-eta2-phi7*/	4, 94, 0, 5, 95, 0, 1, 95, 1, 12, 124, 0, 4, 
/* out0143_had-eta3-phi7*/	9, 64, 2, 1, 93, 0, 14, 93, 2, 7, 94, 0, 4, 94, 1, 1, 95, 0, 10, 95, 1, 4, 123, 0, 1, 124, 0, 4, 
/* out0144_had-eta4-phi7*/	5, 63, 2, 9, 91, 0, 6, 93, 0, 2, 93, 1, 14, 123, 0, 4, 
/* out0145_had-eta5-phi7*/	8, 62, 0, 5, 62, 2, 5, 63, 1, 3, 63, 2, 4, 91, 0, 4, 91, 1, 4, 122, 0, 1, 123, 0, 3, 
/* out0146_had-eta6-phi7*/	4, 62, 0, 3, 62, 1, 11, 62, 2, 7, 122, 0, 3, 
/* out0147_had-eta7-phi7*/	4, 61, 0, 14, 62, 1, 2, 71, 2, 2, 122, 0, 3, 
/* out0148_had-eta8-phi7*/	4, 61, 0, 1, 61, 1, 8, 70, 2, 6, 122, 0, 1, 
/* out0149_had-eta9-phi7*/	3, 60, 0, 1, 70, 1, 2, 70, 2, 9, 
/* out0150_had-eta10-phi7*/	6, 8, 0, 3, 8, 2, 2, 8, 3, 16, 8, 9, 6, 8, 10, 1, 70, 1, 2, 
/* out0151_had-eta11-phi7*/	4, 8, 1, 1, 8, 2, 14, 8, 6, 11, 8, 10, 7, 
/* out0152_had-eta12-phi7*/	6, 7, 0, 1, 8, 4, 14, 8, 5, 3, 8, 6, 4, 8, 7, 5, 10, 8, 1, 
/* out0153_had-eta13-phi7*/	4, 7, 0, 11, 7, 1, 3, 10, 8, 8, 10, 11, 1, 
/* out0154_had-eta14-phi7*/	3, 7, 1, 11, 7, 7, 4, 10, 11, 4, 
/* out0155_had-eta15-phi7*/	3, 7, 7, 3, 9, 3, 1, 9, 9, 12, 
/* out0156_had-eta16-phi7*/	2, 9, 9, 4, 9, 10, 9, 
/* out0157_had-eta17-phi7*/	3, 9, 6, 4, 9, 10, 6, 9, 11, 2, 
/* out0158_had-eta18-phi7*/	1, 9, 5, 9, 
/* out0159_had-eta19-phi7*/	2, 9, 4, 2, 9, 5, 1, 
/* out0160_had-eta0-phi8*/	1, 129, 0, 4, 
/* out0161_had-eta1-phi8*/	1, 129, 0, 4, 
/* out0162_had-eta2-phi8*/	1, 128, 0, 4, 
/* out0163_had-eta3-phi8*/	6, 64, 0, 11, 64, 1, 5, 64, 2, 14, 95, 0, 5, 127, 0, 1, 128, 0, 4, 
/* out0164_had-eta4-phi8*/	6, 63, 0, 15, 63, 2, 3, 64, 1, 9, 64, 2, 1, 73, 2, 3, 127, 0, 4, 
/* out0165_had-eta5-phi8*/	6, 62, 0, 3, 63, 0, 1, 63, 1, 13, 72, 2, 9, 126, 0, 1, 127, 0, 3, 
/* out0166_had-eta6-phi8*/	7, 62, 0, 5, 62, 1, 3, 71, 0, 3, 71, 2, 2, 72, 1, 3, 72, 2, 5, 126, 0, 3, 
/* out0167_had-eta7-phi8*/	4, 71, 0, 3, 71, 1, 3, 71, 2, 11, 126, 0, 3, 
/* out0168_had-eta8-phi8*/	4, 70, 0, 8, 71, 1, 6, 71, 2, 1, 126, 0, 1, 
/* out0169_had-eta9-phi8*/	3, 70, 0, 5, 70, 1, 6, 70, 2, 1, 
/* out0170_had-eta10-phi8*/	3, 8, 0, 9, 11, 8, 13, 70, 1, 5, 
/* out0171_had-eta11-phi8*/	6, 8, 0, 4, 8, 1, 15, 8, 7, 3, 11, 5, 1, 11, 8, 2, 11, 11, 9, 
/* out0172_had-eta12-phi8*/	6, 8, 4, 1, 8, 7, 8, 10, 3, 2, 10, 8, 3, 10, 9, 14, 10, 10, 1, 
/* out0173_had-eta13-phi8*/	4, 10, 8, 4, 10, 9, 2, 10, 10, 12, 10, 11, 5, 
/* out0174_had-eta14-phi8*/	4, 10, 5, 11, 10, 6, 2, 10, 10, 1, 10, 11, 6, 
/* out0175_had-eta15-phi8*/	3, 9, 0, 1, 9, 3, 13, 10, 5, 2, 
/* out0176_had-eta16-phi8*/	3, 9, 2, 11, 9, 3, 2, 9, 10, 1, 
/* out0177_had-eta17-phi8*/	2, 9, 2, 2, 9, 6, 9, 
/* out0178_had-eta18-phi8*/	4, 9, 4, 5, 9, 5, 1, 9, 6, 2, 9, 7, 2, 
/* out0179_had-eta19-phi8*/	1, 9, 4, 5, 
/* out0180_had-eta0-phi9*/	1, 129, 0, 4, 
/* out0181_had-eta1-phi9*/	1, 129, 0, 4, 
/* out0182_had-eta2-phi9*/	3, 74, 0, 3, 74, 2, 1, 128, 0, 4, 
/* out0183_had-eta3-phi9*/	8, 64, 0, 5, 64, 1, 1, 73, 0, 1, 74, 0, 4, 74, 1, 9, 74, 2, 15, 127, 0, 1, 128, 0, 4, 
/* out0184_had-eta4-phi9*/	5, 64, 1, 1, 73, 0, 11, 73, 1, 7, 73, 2, 12, 127, 0, 4, 
/* out0185_had-eta5-phi9*/	7, 72, 0, 15, 72, 2, 2, 73, 1, 7, 73, 2, 1, 82, 2, 2, 126, 0, 1, 127, 0, 3, 
/* out0186_had-eta6-phi9*/	5, 71, 0, 2, 72, 0, 1, 72, 1, 13, 81, 2, 4, 126, 0, 3, 
/* out0187_had-eta7-phi9*/	5, 71, 0, 8, 71, 1, 4, 80, 0, 1, 81, 2, 4, 126, 0, 3, 
/* out0188_had-eta8-phi9*/	4, 70, 0, 1, 71, 1, 3, 80, 2, 11, 126, 0, 1, 
/* out0189_had-eta9-phi9*/	6, 11, 3, 6, 11, 9, 3, 70, 0, 2, 70, 1, 1, 80, 1, 3, 80, 2, 4, 
/* out0190_had-eta10-phi9*/	6, 11, 2, 7, 11, 3, 6, 11, 8, 1, 11, 9, 13, 11, 10, 11, 11, 11, 1, 
/* out0191_had-eta11-phi9*/	5, 11, 4, 1, 11, 5, 12, 11, 6, 9, 11, 10, 5, 11, 11, 6, 
/* out0192_had-eta12-phi9*/	5, 10, 0, 6, 10, 2, 2, 10, 3, 14, 11, 4, 3, 11, 5, 3, 
/* out0193_had-eta13-phi9*/	4, 10, 1, 1, 10, 2, 13, 10, 6, 7, 10, 10, 2, 
/* out0194_had-eta14-phi9*/	4, 10, 4, 6, 10, 5, 3, 10, 6, 7, 10, 7, 3, 
/* out0195_had-eta15-phi9*/	3, 9, 0, 9, 10, 4, 7, 14, 8, 1, 
/* out0196_had-eta16-phi9*/	3, 9, 0, 5, 9, 1, 7, 9, 2, 2, 
/* out0197_had-eta17-phi9*/	4, 9, 1, 4, 9, 2, 1, 9, 6, 1, 9, 7, 5, 
/* out0198_had-eta18-phi9*/	3, 9, 4, 3, 9, 7, 6, 12, 4, 3, 
/* out0199_had-eta19-phi9*/	2, 9, 4, 1, 12, 4, 11, 
/* out0200_had-eta0-phi10*/	1, 133, 0, 4, 
/* out0201_had-eta1-phi10*/	1, 133, 0, 4, 
/* out0202_had-eta2-phi10*/	3, 74, 0, 1, 84, 1, 3, 132, 0, 4, 
/* out0203_had-eta3-phi10*/	8, 74, 0, 8, 74, 1, 7, 83, 0, 6, 83, 2, 6, 84, 0, 6, 84, 1, 13, 131, 0, 1, 132, 0, 4, 
/* out0204_had-eta4-phi10*/	8, 73, 0, 4, 73, 1, 2, 82, 0, 4, 82, 2, 1, 83, 0, 1, 83, 1, 8, 83, 2, 10, 131, 0, 4, 
/* out0205_had-eta5-phi10*/	5, 82, 0, 6, 82, 1, 7, 82, 2, 13, 130, 0, 1, 131, 0, 3, 
/* out0206_had-eta6-phi10*/	4, 81, 0, 11, 81, 2, 5, 82, 1, 4, 130, 0, 3, 
/* out0207_had-eta7-phi10*/	4, 80, 0, 2, 81, 1, 13, 81, 2, 3, 130, 0, 3, 
/* out0208_had-eta8-phi10*/	4, 80, 0, 11, 80, 1, 2, 80, 2, 1, 130, 0, 1, 
/* out0209_had-eta9-phi10*/	4, 11, 0, 4, 11, 3, 1, 28, 2, 1, 80, 1, 10, 
/* out0210_had-eta10-phi10*/	5, 11, 0, 12, 11, 1, 12, 11, 2, 9, 11, 3, 3, 28, 2, 1, 
/* out0211_had-eta11-phi10*/	6, 11, 1, 2, 11, 4, 7, 11, 6, 7, 11, 7, 14, 15, 8, 1, 15, 9, 1, 
/* out0212_had-eta12-phi10*/	4, 10, 0, 9, 11, 4, 5, 15, 8, 13, 15, 11, 1, 
/* out0213_had-eta13-phi10*/	5, 10, 0, 1, 10, 1, 15, 10, 2, 1, 10, 7, 3, 15, 11, 3, 
/* out0214_had-eta14-phi10*/	4, 10, 4, 2, 10, 7, 10, 14, 8, 1, 14, 9, 5, 
/* out0215_had-eta15-phi10*/	4, 10, 4, 1, 14, 8, 12, 14, 9, 2, 14, 11, 1, 
/* out0216_had-eta16-phi10*/	4, 9, 0, 1, 9, 1, 2, 14, 8, 2, 14, 11, 8, 
/* out0217_had-eta17-phi10*/	6, 9, 1, 3, 9, 7, 2, 12, 3, 1, 12, 5, 1, 14, 5, 1, 14, 11, 3, 
/* out0218_had-eta18-phi10*/	2, 9, 7, 1, 12, 5, 9, 
/* out0219_had-eta19-phi10*/	3, 12, 4, 2, 12, 5, 4, 12, 6, 1, 
/* out0220_had-eta0-phi11*/	1, 133, 0, 4, 
/* out0221_had-eta1-phi11*/	1, 133, 0, 4, 
/* out0222_had-eta2-phi11*/	1, 132, 0, 4, 
/* out0223_had-eta3-phi11*/	4, 83, 0, 6, 84, 0, 10, 131, 0, 1, 132, 0, 4, 
/* out0224_had-eta4-phi11*/	6, 31, 0, 4, 31, 2, 11, 82, 0, 1, 83, 0, 3, 83, 1, 8, 131, 0, 4, 
/* out0225_had-eta5-phi11*/	8, 30, 0, 3, 30, 2, 3, 31, 1, 4, 31, 2, 5, 82, 0, 5, 82, 1, 4, 130, 0, 1, 131, 0, 3, 
/* out0226_had-eta6-phi11*/	6, 30, 0, 1, 30, 1, 3, 30, 2, 13, 81, 0, 4, 82, 1, 1, 130, 0, 3, 
/* out0227_had-eta7-phi11*/	6, 29, 0, 4, 29, 2, 9, 30, 1, 1, 81, 0, 1, 81, 1, 3, 130, 0, 3, 
/* out0228_had-eta8-phi11*/	4, 29, 1, 4, 29, 2, 7, 80, 0, 2, 130, 0, 1, 
/* out0229_had-eta9-phi11*/	3, 28, 0, 3, 28, 2, 8, 80, 1, 1, 
/* out0230_had-eta10-phi11*/	3, 11, 1, 1, 28, 1, 3, 28, 2, 6, 
/* out0231_had-eta11-phi11*/	7, 11, 1, 1, 11, 7, 2, 15, 2, 2, 15, 3, 12, 15, 9, 12, 15, 10, 1, 28, 1, 1, 
/* out0232_had-eta12-phi11*/	6, 15, 2, 2, 15, 6, 2, 15, 8, 2, 15, 9, 3, 15, 10, 15, 15, 11, 4, 
/* out0233_had-eta13-phi11*/	4, 14, 3, 1, 15, 5, 12, 15, 6, 2, 15, 11, 8, 
/* out0234_had-eta14-phi11*/	4, 14, 2, 2, 14, 3, 10, 14, 9, 7, 14, 10, 1, 
/* out0235_had-eta15-phi11*/	4, 14, 2, 2, 14, 6, 1, 14, 9, 2, 14, 10, 12, 
/* out0236_had-eta16-phi11*/	4, 14, 5, 3, 14, 6, 3, 14, 10, 3, 14, 11, 4, 
/* out0237_had-eta17-phi11*/	2, 12, 3, 3, 14, 5, 8, 
/* out0238_had-eta18-phi11*/	3, 12, 2, 1, 12, 3, 8, 12, 5, 1, 
/* out0239_had-eta19-phi11*/	3, 12, 2, 4, 12, 5, 1, 12, 6, 15, 
/* out0240_had-eta0-phi12*/	1, 137, 0, 4, 
/* out0241_had-eta1-phi12*/	1, 137, 0, 4, 
/* out0242_had-eta2-phi12*/	1, 136, 0, 4, 
/* out0243_had-eta3-phi12*/	6, 40, 0, 2, 40, 2, 4, 41, 0, 2, 41, 1, 16, 135, 0, 1, 136, 0, 4, 
/* out0244_had-eta4-phi12*/	6, 31, 0, 12, 31, 1, 4, 39, 2, 1, 40, 1, 1, 40, 2, 10, 135, 0, 4, 
/* out0245_had-eta5-phi12*/	5, 30, 0, 7, 31, 1, 8, 39, 2, 10, 134, 0, 1, 135, 0, 3, 
/* out0246_had-eta6-phi12*/	5, 30, 0, 5, 30, 1, 11, 38, 2, 4, 39, 2, 1, 134, 0, 3, 
/* out0247_had-eta7-phi12*/	5, 29, 0, 12, 29, 1, 1, 30, 1, 1, 38, 2, 4, 134, 0, 3, 
/* out0248_had-eta8-phi12*/	4, 28, 0, 1, 29, 1, 11, 37, 2, 2, 134, 0, 1, 
/* out0249_had-eta9-phi12*/	2, 28, 0, 11, 37, 2, 1, 
/* out0250_had-eta10-phi12*/	2, 18, 8, 1, 28, 1, 10, 
/* out0251_had-eta11-phi12*/	6, 15, 0, 15, 15, 1, 4, 15, 2, 3, 15, 3, 4, 18, 8, 3, 28, 1, 1, 
/* out0252_had-eta12-phi12*/	4, 15, 1, 4, 15, 2, 9, 15, 6, 10, 15, 7, 5, 
/* out0253_had-eta13-phi12*/	5, 14, 0, 1, 15, 4, 13, 15, 5, 4, 15, 6, 2, 15, 7, 2, 
/* out0254_had-eta14-phi12*/	4, 14, 0, 11, 14, 1, 2, 14, 2, 2, 14, 3, 5, 
/* out0255_had-eta15-phi12*/	3, 14, 1, 1, 14, 2, 10, 14, 6, 5, 
/* out0256_had-eta16-phi12*/	4, 14, 4, 2, 14, 5, 2, 14, 6, 7, 14, 7, 2, 
/* out0257_had-eta17-phi12*/	3, 12, 0, 3, 14, 4, 6, 14, 5, 2, 
/* out0258_had-eta18-phi12*/	3, 12, 0, 4, 12, 2, 1, 12, 3, 4, 
/* out0259_had-eta19-phi12*/	1, 12, 2, 9, 
/* out0260_had-eta0-phi13*/	1, 137, 0, 4, 
/* out0261_had-eta1-phi13*/	1, 137, 0, 4, 
/* out0262_had-eta2-phi13*/	3, 41, 0, 2, 51, 0, 1, 136, 0, 4, 
/* out0263_had-eta3-phi13*/	6, 40, 0, 11, 41, 0, 12, 51, 0, 1, 51, 2, 14, 135, 0, 1, 136, 0, 4, 
/* out0264_had-eta4-phi13*/	6, 39, 0, 5, 40, 0, 3, 40, 1, 15, 40, 2, 2, 50, 2, 6, 135, 0, 4, 
/* out0265_had-eta5-phi13*/	5, 39, 0, 10, 39, 1, 11, 39, 2, 4, 134, 0, 1, 135, 0, 3, 
/* out0266_had-eta6-phi13*/	4, 38, 0, 13, 38, 2, 3, 39, 1, 4, 134, 0, 3, 
/* out0267_had-eta7-phi13*/	4, 37, 0, 2, 38, 1, 10, 38, 2, 5, 134, 0, 3, 
/* out0268_had-eta8-phi13*/	4, 37, 0, 6, 37, 1, 1, 37, 2, 8, 134, 0, 1, 
/* out0269_had-eta9-phi13*/	4, 18, 3, 4, 28, 0, 1, 37, 1, 5, 37, 2, 5, 
/* out0270_had-eta10-phi13*/	6, 18, 2, 2, 18, 3, 8, 18, 8, 4, 18, 9, 16, 18, 10, 7, 28, 1, 1, 
/* out0271_had-eta11-phi13*/	6, 15, 0, 1, 15, 1, 2, 18, 5, 2, 18, 8, 8, 18, 10, 7, 18, 11, 14, 
/* out0272_had-eta12-phi13*/	6, 15, 1, 6, 15, 7, 8, 16, 3, 2, 16, 9, 6, 18, 5, 3, 18, 11, 2, 
/* out0273_had-eta13-phi13*/	5, 15, 4, 3, 15, 7, 1, 16, 8, 11, 16, 9, 8, 16, 10, 1, 
/* out0274_had-eta14-phi13*/	4, 14, 0, 4, 14, 1, 4, 16, 8, 5, 16, 11, 7, 
/* out0275_had-eta15-phi13*/	2, 14, 1, 9, 14, 7, 6, 
/* out0276_had-eta16-phi13*/	4, 13, 8, 2, 13, 9, 1, 14, 4, 4, 14, 7, 7, 
/* out0277_had-eta17-phi13*/	3, 12, 0, 2, 13, 8, 6, 14, 4, 4, 
/* out0278_had-eta18-phi13*/	3, 12, 0, 7, 12, 1, 3, 13, 8, 1, 
/* out0279_had-eta19-phi13*/	2, 12, 1, 7, 12, 2, 1, 
/* out0280_had-eta0-phi14*/	1, 141, 0, 4, 
/* out0281_had-eta1-phi14*/	1, 141, 0, 4, 
/* out0282_had-eta2-phi14*/	2, 51, 0, 4, 140, 0, 4, 
/* out0283_had-eta3-phi14*/	7, 50, 0, 1, 51, 0, 10, 51, 1, 16, 51, 2, 2, 59, 2, 6, 139, 0, 1, 140, 0, 4, 
/* out0284_had-eta4-phi14*/	5, 50, 0, 14, 50, 1, 9, 50, 2, 8, 59, 2, 1, 139, 0, 4, 
/* out0285_had-eta5-phi14*/	8, 39, 0, 1, 39, 1, 1, 49, 0, 10, 49, 2, 7, 50, 1, 5, 50, 2, 2, 138, 0, 1, 139, 0, 3, 
/* out0286_had-eta6-phi14*/	6, 38, 0, 3, 38, 1, 1, 48, 0, 2, 49, 1, 6, 49, 2, 9, 138, 0, 3, 
/* out0287_had-eta7-phi14*/	5, 37, 0, 1, 38, 1, 5, 48, 0, 1, 48, 2, 11, 138, 0, 3, 
/* out0288_had-eta8-phi14*/	5, 37, 0, 7, 37, 1, 4, 47, 2, 1, 48, 2, 3, 138, 0, 1, 
/* out0289_had-eta9-phi14*/	3, 18, 0, 8, 37, 1, 6, 47, 2, 3, 
/* out0290_had-eta10-phi14*/	7, 18, 0, 8, 18, 1, 9, 18, 2, 14, 18, 3, 4, 18, 6, 3, 18, 7, 1, 18, 10, 1, 
/* out0291_had-eta11-phi14*/	5, 18, 4, 7, 18, 5, 8, 18, 6, 13, 18, 7, 4, 18, 10, 1, 
/* out0292_had-eta12-phi14*/	6, 16, 0, 6, 16, 2, 2, 16, 3, 14, 16, 9, 1, 18, 4, 2, 18, 5, 3, 
/* out0293_had-eta13-phi14*/	4, 16, 2, 8, 16, 6, 2, 16, 9, 1, 16, 10, 12, 
/* out0294_had-eta14-phi14*/	4, 16, 5, 6, 16, 6, 4, 16, 10, 3, 16, 11, 7, 
/* out0295_had-eta15-phi14*/	5, 13, 3, 6, 13, 9, 3, 14, 7, 1, 16, 5, 5, 16, 11, 2, 
/* out0296_had-eta16-phi14*/	3, 13, 3, 1, 13, 9, 11, 13, 10, 1, 
/* out0297_had-eta17-phi14*/	4, 13, 8, 5, 13, 9, 1, 13, 10, 3, 13, 11, 2, 
/* out0298_had-eta18-phi14*/	3, 12, 1, 2, 13, 8, 2, 13, 11, 7, 
/* out0299_had-eta19-phi14*/	2, 12, 1, 4, 13, 11, 1, 
/* out0300_had-eta0-phi15*/	1, 141, 0, 4, 
/* out0301_had-eta1-phi15*/	1, 141, 0, 4, 
/* out0302_had-eta2-phi15*/	1, 140, 0, 4, 
/* out0303_had-eta3-phi15*/	6, 59, 0, 16, 59, 1, 8, 59, 2, 6, 109, 1, 9, 139, 0, 1, 140, 0, 4, 
/* out0304_had-eta4-phi15*/	7, 50, 0, 1, 50, 1, 2, 58, 0, 10, 58, 2, 7, 59, 1, 7, 59, 2, 3, 139, 0, 4, 
/* out0305_had-eta5-phi15*/	8, 49, 0, 6, 49, 1, 3, 57, 0, 2, 57, 2, 1, 58, 1, 5, 58, 2, 9, 138, 0, 1, 139, 0, 3, 
/* out0306_had-eta6-phi15*/	4, 48, 0, 5, 49, 1, 7, 57, 2, 9, 138, 0, 3, 
/* out0307_had-eta7-phi15*/	4, 48, 0, 8, 48, 1, 8, 48, 2, 2, 138, 0, 3, 
/* out0308_had-eta8-phi15*/	4, 47, 0, 7, 47, 2, 1, 48, 1, 6, 138, 0, 1, 
/* out0309_had-eta9-phi15*/	3, 47, 0, 2, 47, 1, 2, 47, 2, 8, 
/* out0310_had-eta10-phi15*/	6, 17, 3, 5, 17, 9, 4, 18, 1, 7, 18, 7, 6, 47, 1, 2, 47, 2, 3, 
/* out0311_had-eta11-phi15*/	4, 17, 8, 10, 17, 9, 11, 18, 4, 7, 18, 7, 5, 
/* out0312_had-eta12-phi15*/	5, 16, 0, 10, 16, 1, 8, 16, 2, 1, 17, 8, 6, 17, 11, 3, 
/* out0313_had-eta13-phi15*/	4, 16, 1, 5, 16, 2, 5, 16, 6, 7, 16, 7, 7, 
/* out0314_had-eta14-phi15*/	4, 16, 4, 10, 16, 5, 4, 16, 6, 3, 16, 7, 2, 
/* out0315_had-eta15-phi15*/	4, 13, 0, 6, 13, 3, 7, 16, 4, 1, 16, 5, 1, 
/* out0316_had-eta16-phi15*/	3, 13, 2, 9, 13, 3, 2, 13, 10, 3, 
/* out0317_had-eta17-phi15*/	2, 13, 6, 3, 13, 10, 8, 
/* out0318_had-eta18-phi15*/	4, 13, 5, 4, 13, 6, 1, 13, 10, 1, 13, 11, 4, 
/* out0319_had-eta19-phi15*/	2, 13, 5, 4, 13, 11, 2, 
/* out0320_had-eta0-phi16*/	1, 145, 0, 4, 
/* out0321_had-eta1-phi16*/	1, 145, 0, 4, 
/* out0322_had-eta2-phi16*/	4, 108, 1, 3, 109, 0, 6, 109, 1, 2, 144, 0, 4, 
/* out0323_had-eta3-phi16*/	9, 59, 1, 1, 107, 0, 14, 107, 1, 2, 107, 2, 7, 108, 1, 3, 109, 0, 10, 109, 1, 5, 143, 0, 1, 144, 0, 4, 
/* out0324_had-eta4-phi16*/	7, 58, 0, 6, 58, 1, 4, 106, 0, 3, 106, 2, 3, 107, 1, 7, 107, 2, 9, 143, 0, 4, 
/* out0325_had-eta5-phi16*/	5, 57, 0, 10, 58, 1, 7, 106, 2, 8, 142, 0, 1, 143, 0, 3, 
/* out0326_had-eta6-phi16*/	4, 57, 0, 4, 57, 1, 12, 57, 2, 5, 142, 0, 3, 
/* out0327_had-eta7-phi16*/	6, 48, 1, 2, 56, 0, 6, 56, 2, 8, 57, 1, 1, 57, 2, 1, 142, 0, 3, 
/* out0328_had-eta8-phi16*/	3, 47, 0, 6, 56, 2, 8, 142, 0, 1, 
/* out0329_had-eta9-phi16*/	3, 47, 0, 1, 47, 1, 9, 65, 2, 1, 
/* out0330_had-eta10-phi16*/	5, 17, 0, 13, 17, 1, 2, 17, 2, 3, 17, 3, 11, 47, 1, 3, 
/* out0331_had-eta11-phi16*/	5, 17, 2, 11, 17, 6, 7, 17, 9, 1, 17, 10, 14, 17, 11, 1, 
/* out0332_had-eta12-phi16*/	5, 16, 1, 1, 17, 5, 10, 17, 6, 2, 17, 10, 2, 17, 11, 12, 
/* out0333_had-eta13-phi16*/	4, 16, 1, 2, 16, 7, 7, 19, 3, 3, 19, 9, 9, 
/* out0334_had-eta14-phi16*/	3, 16, 4, 5, 19, 8, 11, 19, 9, 2, 
/* out0335_had-eta15-phi16*/	3, 13, 0, 10, 13, 1, 4, 19, 8, 2, 
/* out0336_had-eta16-phi16*/	3, 13, 1, 4, 13, 2, 7, 13, 6, 2, 
/* out0337_had-eta17-phi16*/	2, 13, 6, 9, 13, 7, 2, 
/* out0338_had-eta18-phi16*/	3, 13, 4, 3, 13, 5, 6, 13, 6, 1, 
/* out0339_had-eta19-phi16*/	1, 13, 5, 2, 
/* out0340_had-eta0-phi17*/	1, 145, 0, 4, 
/* out0341_had-eta1-phi17*/	1, 145, 0, 4, 
/* out0342_had-eta2-phi17*/	2, 108, 1, 2, 144, 0, 4, 
/* out0343_had-eta3-phi17*/	8, 100, 0, 8, 100, 2, 4, 107, 0, 2, 107, 1, 3, 108, 0, 16, 108, 1, 8, 143, 0, 1, 144, 0, 4, 
/* out0344_had-eta4-phi17*/	5, 100, 2, 12, 106, 0, 12, 106, 1, 2, 107, 1, 4, 143, 0, 4, 
/* out0345_had-eta5-phi17*/	6, 96, 0, 5, 106, 0, 1, 106, 1, 14, 106, 2, 5, 142, 0, 1, 143, 0, 3, 
/* out0346_had-eta6-phi17*/	5, 56, 0, 1, 57, 1, 3, 96, 0, 3, 96, 2, 14, 142, 0, 3, 
/* out0347_had-eta7-phi17*/	4, 56, 0, 9, 56, 1, 7, 96, 2, 2, 142, 0, 3, 
/* out0348_had-eta8-phi17*/	3, 56, 1, 9, 65, 0, 4, 142, 0, 1, 
/* out0349_had-eta9-phi17*/	2, 65, 0, 3, 65, 2, 9, 
/* out0350_had-eta10-phi17*/	4, 17, 0, 3, 17, 1, 12, 17, 7, 1, 65, 2, 6, 
/* out0351_had-eta11-phi17*/	5, 17, 1, 2, 17, 2, 2, 17, 4, 5, 17, 6, 7, 17, 7, 15, 
/* out0352_had-eta12-phi17*/	4, 17, 4, 11, 17, 5, 6, 19, 0, 7, 19, 3, 3, 
/* out0353_had-eta13-phi17*/	4, 19, 2, 7, 19, 3, 10, 19, 9, 3, 19, 10, 3, 
/* out0354_had-eta14-phi17*/	4, 19, 8, 2, 19, 9, 2, 19, 10, 12, 19, 11, 3, 
/* out0355_had-eta15-phi17*/	3, 13, 1, 3, 19, 8, 1, 19, 11, 12, 
/* out0356_had-eta16-phi17*/	2, 13, 1, 5, 13, 7, 8, 
/* out0357_had-eta17-phi17*/	2, 13, 4, 5, 13, 7, 6, 
/* out0358_had-eta18-phi17*/	1, 13, 4, 8, 
/* out0359_had-eta19-phi17*/	0, 
/* out0360_had-eta0-phi18*/	1, 149, 0, 4, 
/* out0361_had-eta1-phi18*/	1, 149, 0, 4, 
/* out0362_had-eta2-phi18*/	2, 101, 0, 2, 148, 0, 4, 
/* out0363_had-eta3-phi18*/	8, 98, 0, 2, 98, 2, 3, 100, 0, 8, 100, 1, 4, 101, 0, 8, 101, 1, 16, 147, 0, 1, 148, 0, 4, 
/* out0364_had-eta4-phi18*/	5, 97, 0, 12, 97, 2, 2, 98, 2, 4, 100, 1, 12, 147, 0, 4, 
/* out0365_had-eta5-phi18*/	6, 96, 0, 5, 97, 0, 1, 97, 1, 5, 97, 2, 14, 146, 0, 1, 147, 0, 3, 
/* out0366_had-eta6-phi18*/	5, 66, 0, 1, 67, 2, 3, 96, 0, 3, 96, 1, 14, 146, 0, 3, 
/* out0367_had-eta7-phi18*/	4, 66, 0, 9, 66, 2, 7, 96, 1, 2, 146, 0, 3, 
/* out0368_had-eta8-phi18*/	3, 65, 0, 5, 66, 2, 9, 146, 0, 1, 
/* out0369_had-eta9-phi18*/	2, 65, 0, 4, 65, 1, 9, 
/* out0370_had-eta10-phi18*/	4, 20, 0, 3, 20, 3, 12, 20, 9, 1, 65, 1, 6, 
/* out0371_had-eta11-phi18*/	5, 20, 2, 2, 20, 3, 2, 20, 8, 5, 20, 9, 15, 20, 10, 7, 
/* out0372_had-eta12-phi18*/	4, 19, 0, 8, 19, 1, 3, 20, 8, 11, 20, 11, 6, 
/* out0373_had-eta13-phi18*/	5, 19, 0, 1, 19, 1, 9, 19, 2, 9, 19, 6, 3, 19, 7, 2, 
/* out0374_had-eta14-phi18*/	5, 19, 4, 1, 19, 5, 4, 19, 6, 13, 19, 7, 1, 19, 10, 1, 
/* out0375_had-eta15-phi18*/	3, 19, 5, 12, 19, 11, 1, 21, 3, 3, 
/* out0376_had-eta16-phi18*/	2, 21, 3, 5, 21, 9, 8, 
/* out0377_had-eta17-phi18*/	2, 21, 8, 5, 21, 9, 6, 
/* out0378_had-eta18-phi18*/	1, 21, 8, 8, 
/* out0379_had-eta19-phi18*/	0, 
/* out0380_had-eta0-phi19*/	1, 149, 0, 4, 
/* out0381_had-eta1-phi19*/	1, 149, 0, 4, 
/* out0382_had-eta2-phi19*/	4, 99, 0, 2, 99, 1, 6, 101, 0, 3, 148, 0, 4, 
/* out0383_had-eta3-phi19*/	9, 69, 2, 1, 98, 0, 14, 98, 1, 7, 98, 2, 2, 99, 0, 5, 99, 1, 10, 101, 0, 3, 147, 0, 1, 148, 0, 4, 
/* out0384_had-eta4-phi19*/	7, 68, 0, 6, 68, 2, 4, 97, 0, 3, 97, 1, 3, 98, 1, 9, 98, 2, 7, 147, 0, 4, 
/* out0385_had-eta5-phi19*/	5, 67, 0, 10, 68, 2, 7, 97, 1, 8, 146, 0, 1, 147, 0, 3, 
/* out0386_had-eta6-phi19*/	4, 67, 0, 4, 67, 1, 5, 67, 2, 12, 146, 0, 3, 
/* out0387_had-eta7-phi19*/	6, 66, 0, 6, 66, 1, 8, 67, 1, 1, 67, 2, 1, 76, 2, 2, 146, 0, 3, 
/* out0388_had-eta8-phi19*/	3, 66, 1, 8, 75, 0, 6, 146, 0, 1, 
/* out0389_had-eta9-phi19*/	3, 65, 1, 1, 75, 0, 1, 75, 2, 9, 
/* out0390_had-eta10-phi19*/	5, 20, 0, 13, 20, 1, 11, 20, 2, 3, 20, 3, 2, 75, 2, 3, 
/* out0391_had-eta11-phi19*/	5, 20, 2, 11, 20, 5, 1, 20, 6, 14, 20, 7, 1, 20, 10, 7, 
/* out0392_had-eta12-phi19*/	6, 19, 1, 1, 20, 5, 12, 20, 6, 2, 20, 10, 2, 20, 11, 10, 22, 3, 1, 
/* out0393_had-eta13-phi19*/	4, 19, 1, 3, 19, 7, 10, 22, 3, 2, 22, 9, 7, 
/* out0394_had-eta14-phi19*/	3, 19, 4, 12, 19, 7, 3, 22, 8, 5, 
/* out0395_had-eta15-phi19*/	3, 19, 4, 3, 21, 0, 10, 21, 3, 4, 
/* out0396_had-eta16-phi19*/	3, 21, 2, 7, 21, 3, 4, 21, 10, 2, 
/* out0397_had-eta17-phi19*/	2, 21, 9, 2, 21, 10, 9, 
/* out0398_had-eta18-phi19*/	3, 21, 8, 3, 21, 10, 1, 21, 11, 6, 
/* out0399_had-eta19-phi19*/	1, 21, 11, 2, 
/* out0400_had-eta0-phi20*/	1, 153, 0, 4, 
/* out0401_had-eta1-phi20*/	1, 153, 0, 4, 
/* out0402_had-eta2-phi20*/	1, 152, 0, 4, 
/* out0403_had-eta3-phi20*/	6, 69, 0, 16, 69, 1, 6, 69, 2, 8, 99, 0, 9, 151, 0, 1, 152, 0, 4, 
/* out0404_had-eta4-phi20*/	7, 68, 0, 10, 68, 1, 7, 69, 1, 3, 69, 2, 7, 78, 0, 1, 78, 2, 2, 151, 0, 4, 
/* out0405_had-eta5-phi20*/	8, 67, 0, 2, 67, 1, 1, 68, 1, 9, 68, 2, 5, 77, 0, 6, 77, 2, 3, 150, 0, 1, 151, 0, 3, 
/* out0406_had-eta6-phi20*/	4, 67, 1, 9, 76, 0, 5, 77, 2, 7, 150, 0, 3, 
/* out0407_had-eta7-phi20*/	4, 76, 0, 8, 76, 1, 2, 76, 2, 8, 150, 0, 3, 
/* out0408_had-eta8-phi20*/	4, 75, 0, 7, 75, 1, 1, 76, 2, 6, 150, 0, 1, 
/* out0409_had-eta9-phi20*/	3, 75, 0, 2, 75, 1, 8, 75, 2, 2, 
/* out0410_had-eta10-phi20*/	6, 20, 1, 5, 20, 7, 4, 23, 3, 7, 23, 9, 6, 75, 1, 3, 75, 2, 2, 
/* out0411_had-eta11-phi20*/	4, 20, 4, 10, 20, 7, 11, 23, 8, 7, 23, 9, 5, 
/* out0412_had-eta12-phi20*/	5, 20, 4, 6, 20, 5, 3, 22, 0, 10, 22, 2, 1, 22, 3, 8, 
/* out0413_had-eta13-phi20*/	4, 22, 2, 5, 22, 3, 5, 22, 9, 7, 22, 10, 7, 
/* out0414_had-eta14-phi20*/	4, 22, 8, 10, 22, 9, 2, 22, 10, 3, 22, 11, 4, 
/* out0415_had-eta15-phi20*/	4, 21, 0, 6, 21, 1, 7, 22, 8, 1, 22, 11, 1, 
/* out0416_had-eta16-phi20*/	3, 21, 1, 2, 21, 2, 9, 21, 6, 3, 
/* out0417_had-eta17-phi20*/	2, 21, 6, 8, 21, 10, 3, 
/* out0418_had-eta18-phi20*/	4, 21, 5, 4, 21, 6, 1, 21, 10, 1, 21, 11, 4, 
/* out0419_had-eta19-phi20*/	2, 21, 5, 2, 21, 11, 4, 
/* out0420_had-eta0-phi21*/	1, 153, 0, 4, 
/* out0421_had-eta1-phi21*/	1, 153, 0, 4, 
/* out0422_had-eta2-phi21*/	2, 79, 0, 4, 152, 0, 4, 
/* out0423_had-eta3-phi21*/	7, 69, 1, 6, 78, 0, 1, 79, 0, 10, 79, 1, 2, 79, 2, 16, 151, 0, 1, 152, 0, 4, 
/* out0424_had-eta4-phi21*/	5, 69, 1, 1, 78, 0, 14, 78, 1, 8, 78, 2, 9, 151, 0, 4, 
/* out0425_had-eta5-phi21*/	8, 77, 0, 10, 77, 1, 7, 78, 1, 2, 78, 2, 5, 87, 0, 1, 87, 2, 1, 150, 0, 1, 151, 0, 3, 
/* out0426_had-eta6-phi21*/	6, 76, 0, 2, 77, 1, 9, 77, 2, 6, 86, 0, 3, 86, 2, 1, 150, 0, 3, 
/* out0427_had-eta7-phi21*/	5, 76, 0, 1, 76, 1, 11, 85, 0, 1, 86, 2, 5, 150, 0, 3, 
/* out0428_had-eta8-phi21*/	5, 75, 1, 1, 76, 1, 3, 85, 0, 7, 85, 2, 4, 150, 0, 1, 
/* out0429_had-eta9-phi21*/	3, 23, 0, 8, 75, 1, 3, 85, 2, 6, 
/* out0430_had-eta10-phi21*/	7, 23, 0, 8, 23, 1, 4, 23, 2, 14, 23, 3, 9, 23, 6, 1, 23, 9, 1, 23, 10, 3, 
/* out0431_had-eta11-phi21*/	5, 23, 6, 1, 23, 8, 7, 23, 9, 4, 23, 10, 13, 23, 11, 8, 
/* out0432_had-eta12-phi21*/	6, 22, 0, 6, 22, 1, 14, 22, 2, 2, 22, 7, 1, 23, 8, 2, 23, 11, 3, 
/* out0433_had-eta13-phi21*/	4, 22, 2, 8, 22, 6, 12, 22, 7, 1, 22, 10, 2, 
/* out0434_had-eta14-phi21*/	4, 22, 5, 7, 22, 6, 3, 22, 10, 4, 22, 11, 6, 
/* out0435_had-eta15-phi21*/	4, 21, 1, 6, 21, 7, 3, 22, 5, 2, 22, 11, 5, 
/* out0436_had-eta16-phi21*/	3, 21, 1, 1, 21, 6, 1, 21, 7, 11, 
/* out0437_had-eta17-phi21*/	4, 21, 4, 5, 21, 5, 2, 21, 6, 3, 21, 7, 1, 
/* out0438_had-eta18-phi21*/	2, 21, 4, 2, 21, 5, 7, 
/* out0439_had-eta19-phi21*/	1, 21, 5, 1, 
/* out0440_had-eta0-phi22*/	1, 157, 0, 4, 
/* out0441_had-eta1-phi22*/	1, 157, 0, 4, 
/* out0442_had-eta2-phi22*/	3, 79, 0, 1, 89, 1, 2, 156, 0, 4, 
/* out0443_had-eta3-phi22*/	6, 79, 0, 1, 79, 1, 14, 88, 0, 11, 89, 1, 12, 155, 0, 1, 156, 0, 4, 
/* out0444_had-eta4-phi22*/	6, 78, 1, 6, 87, 0, 5, 88, 0, 3, 88, 1, 2, 88, 2, 15, 155, 0, 4, 
/* out0445_had-eta5-phi22*/	5, 87, 0, 10, 87, 1, 4, 87, 2, 11, 154, 0, 1, 155, 0, 3, 
/* out0446_had-eta6-phi22*/	4, 86, 0, 13, 86, 1, 3, 87, 2, 4, 154, 0, 3, 
/* out0447_had-eta7-phi22*/	4, 85, 0, 2, 86, 1, 5, 86, 2, 10, 154, 0, 3, 
/* out0448_had-eta8-phi22*/	4, 85, 0, 6, 85, 1, 8, 85, 2, 1, 154, 0, 1, 
/* out0449_had-eta9-phi22*/	3, 23, 1, 4, 85, 1, 5, 85, 2, 5, 
/* out0450_had-eta10-phi22*/	5, 23, 1, 8, 23, 2, 2, 23, 4, 4, 23, 6, 7, 23, 7, 16, 
/* out0451_had-eta11-phi22*/	4, 23, 4, 8, 23, 5, 14, 23, 6, 7, 23, 11, 2, 
/* out0452_had-eta12-phi22*/	4, 22, 1, 2, 22, 7, 6, 23, 5, 2, 23, 11, 3, 
/* out0453_had-eta13-phi22*/	3, 22, 4, 11, 22, 6, 1, 22, 7, 8, 
/* out0454_had-eta14-phi22*/	2, 22, 4, 5, 22, 5, 7, 
/* out0455_had-eta15-phi22*/	0, 
/* out0456_had-eta16-phi22*/	2, 21, 4, 2, 21, 7, 1, 
/* out0457_had-eta17-phi22*/	1, 21, 4, 6, 
/* out0458_had-eta18-phi22*/	1, 21, 4, 1, 
/* out0459_had-eta19-phi22*/	0, 
/* out0460_had-eta0-phi23*/	1, 157, 0, 4, 
/* out0461_had-eta1-phi23*/	1, 157, 0, 4, 
/* out0462_had-eta2-phi23*/	1, 156, 0, 4, 
/* out0463_had-eta3-phi23*/	6, 88, 0, 2, 88, 1, 4, 89, 0, 16, 89, 1, 2, 155, 0, 1, 156, 0, 4, 
/* out0464_had-eta4-phi23*/	4, 87, 1, 1, 88, 1, 10, 88, 2, 1, 155, 0, 4, 
/* out0465_had-eta5-phi23*/	3, 87, 1, 10, 154, 0, 1, 155, 0, 3, 
/* out0466_had-eta6-phi23*/	3, 86, 1, 4, 87, 1, 1, 154, 0, 3, 
/* out0467_had-eta7-phi23*/	2, 86, 1, 4, 154, 0, 3, 
/* out0468_had-eta8-phi23*/	2, 85, 1, 2, 154, 0, 1, 
/* out0469_had-eta9-phi23*/	1, 85, 1, 1, 
/* out0470_had-eta10-phi23*/	1, 23, 4, 1, 
/* out0471_had-eta11-phi23*/	1, 23, 4, 3, 
/* out0472_had-eta12-phi23*/	0, 
/* out0473_had-eta13-phi23*/	0, 
/* out0474_had-eta14-phi23*/	0, 
/* out0475_had-eta15-phi23*/	0, 
/* out0476_had-eta16-phi23*/	0, 
/* out0477_had-eta17-phi23*/	0, 
/* out0478_had-eta18-phi23*/	0, 
/* out0479_had-eta19-phi23*/	0, 
};